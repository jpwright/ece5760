��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F��T3�y��xq)��8�<LS�A��{Cr��0:���sq��l9���<gJs*UjV����|*���	�k2$�2y���IsM���Ӕ�rJ�2Ɠ�T���ǹ�[�tzR�Фu��@:V\���
p_����%q'Y۴C+H��IDi�ި����.�S/� w����
ٙ�Rp�̕t;�D����M�yބ�{=��;"�*��V��qX��퍶R��E�v2�[y<鵅�,�#��fy'_I�s/�Aݤ�ʫN �M�*K
�u��R�,��L"�����-f�S��������Θb��a�a4p�$d��U�N�ɮ�$��XS��?Px��/�d�E��4��V&K�I ��h(�[>�h<�ջL$�q�;p� lx�ؼ�|�q)�lO$�H�s��u=�_|���0����@�t8�I,�ol��/�]�n+�����4��g6�HҏE��f2�~��)59�:���K�cc�s��&�L���6ϝF������/_� @��pGi��m�����rv`�KطR_��4�~D���AO*�X���4������x����)S]��v�/��=�h��6�;�|U`�FO+�1�dB h�I�PN��(0Z�?�H:��5�i��8��g���6	��|�埫+N@�X{"��e���RhI��M���	�&�d.�s�W�ፖ����>����91L*Ҹ\ A���r��f��a#Ȳ*��F(��;�u��٬JO�0���{kqzpY�����}0R�`��2���,�ҌR�7P�'_��M�+�3P˫}�ژ��|�܀F:��ͣ?8�@�S��
�!7���a���I����%R�n����IQ]9�	˙;�Ӳ�;�x�����h��0܄�Y~��s��E`3`*V /�?*;X��O{�sp� �1n�G/hN>��q-�qZCT�3F%{#Gt*�k�᣼פ�rE� L<&{��'�FքJq��������i�b�|���_#���P��,N,��V-�	�y*y!*
����vɺ����㏣fEM��+
��O)���~���X#ޛ��hm��c�{� �	Wa����4ɍGhg���~�i 1EPvD�LFC��/�O�§X�	���]��?Y�Ȕ	�=� �5�:x�]��k���8K,�㗭�;�yaI{o-r�*-��h�M� �^���Yx��jk��K||`��	�K\��oB��:��M,������w-iG�$b�:�F����>*j�d����K����v�V��"��O�0X�3�e������z���j�\�.�S�M��h�UF��8���hz��TW���;��V��O�8��g��3Hi�l��)q8u�78��ɗ�9Xی�8N��/m~����h���u|�%�����Т�맆�sS�NzQ�� $��DwJ&N��ą��טU9��.�^�/K��ڢc=��3���7I����A�6�miya�֦��f�rςQ(B�q��� p�/�U������.�A�e�lv�B�y_.K���$�<�eX
 
=�����;q~���,y����)To*���!��OUS��).���,C�bV�5�v��T�[�o�<s�UZ؆�5
Z�����V6|@��.�
�^:e
�j�C)�Z���6��E�����s����E���˅�m�#&���	=,��YAD�M�A���t,���t�����X�M�L��S%��iQw0��VǬM�)r�s�{���VZ��)Z���1�'���yת�#����u��L�N
qu��Y.Ւx���Y������Xu��|��������"c��f�1�=m���y�����|�τr����YHd�(?��7`#�����R@j1���=
hm��J=l�����$ٮ���E|�i�l:��2~���i��S��ܧ��bn��k`���ґ"���m<(͜�NN��&�!t�EVwl:�%�V$71d��a�3މ^����t*�(/Tl}XYH�a8��?������n=�ZR���j�	�=|�뒱���B(���͜��َf�"�k���Y���6zk2z�,����w���³V�KXJ-|N�'�2���?w63o��	()Ǡ�M1j������c�-6i>�F+���%��yq�RvK_.yKI�-�7<S�[S��1��t�ύu(�*|m�{���>v���~%�Q=wO��a=�H_�6#�d�^����� ��o&���֐�#Ԋ������_`?�$�r��m A����8�Ӌ'�U%�1��%�N��,��s�p�Pkym�AEXHB��Gm��V+��A��K���ke�_8M��_�
��|W�Q���(�`�I�\���}��
��t�E�7�u�Am�]��ښ6�/���|�6�����}^���'�M�Sz��[�o��xv���M�{xvӊ�ڨkL�>s�5���Ta_B��#['�CsvU����8�a��	�^+�yܖ���]UwT�rqLju�ݳm��c�P��9�\R^��	l�wZ��SY�O�W"�� �U���ko9��4����c��v�nJg�f�J���������̇'w�?,)��n�ذM�G1�Po���s�	�6��m��֌oة�L��n*)�l�mm#��q�'K��E���ܷ���{�M��9��`Ҹ]!�f+�a��`�S*^��qujò������ܖn�#���叭�n�&U�~�r����w�-���p: ���+��4D���@��z!��1ޘ�N	��M��[��/�܈N������E�P�*�Ï2�ʙr��=�C#t��p�W3�^F�k 
R��:���l�U�_���������1�o�m��U/�teI ��pXT!��N�j��[�✎#k���u7D�ڇ�r���gQT���Rը3�J�)su���l$��Km)�=ޠ7�N�@E�����
�����Y)�ϻ������c���]�q��0��\[i��]�Z ��ylh�ȡ-�*��H�Ỵ*~;���)���,H���ڝc��S�ۥ#-�	V+>�Pd� ��tq��Ki�'U:K�y� � W�����|?��ѭ¥��K���t�a�j��;ނ��E����m���4jX<����տ���ک\}���PM�1g�[s��~�B�O���Y7����o�q�΄�f�d�-�R��Q�a`������½hX�t-�wvc��PԜ%T�e�O]���Һ���/Ho�{����F>��Ӥ��&�|��9z=�=�X����
+�:������6�Ky���f{�է�3LQ��W9��T��P�G雪"�;o Fr	�oK�1����l������_��r���[;�`C��'���'�VqzF�vU�/Q�I9 ���y�*䏞�HAʼ���4����F	D�a���"b��!��|&6�'���z�Ά�̶��ďJ]��9V6�P�����Ѿ�9j�(���]�	*���q��݈+��;�2 �h>�8��=�]�Zs_��Y���;��(lP��	���{y�P4JTW��6�6"��������x��H�Cڳ�[�{+�kz�?B�4y�����I��m���:d}�'q>�XYLv����4�������Cj�Z*����naWg/"���b)� ��,�zlS3W��l��y�fa=��A�O�V�#9p9LХ�C�	Q�LB0.oS�,�^/b9�6��n�CP:_��3��X7��7�9Q!K1$���0���*�PK`��Xw����;�f)Zv����n�T[�z�cDF��z90䠝�M�V[�{�(ˡ�����AA��O�A�ɕ���+1��qd4D��۾h�pVB#h�{&���*��{��ܼgi����2��5��D�L��w�w\]��e	�Al#��~U��҃�Fp)��a�g��A���.�]����$c��̏ .�]�!=Ǜz�m.sZ��r�`�1�MU��jz�x+T~=�G�3p|m݅���e�l���'�$������
A���i�[
�s��hy1����O-�?�� �ͺ��"��gM6-����� ��_�^LX�~fI��iǵ
ɐ��͝'&`ʆg(��N�4X妎N��2�C$_�����)e���U���Ki7&��M|V��B�R���n�w䙿���l���A�k,BV��EEF�ƪ��|��<���bCk^�����xԱ����!���Ϩ1-Wv�b]Ǌ�P�>��$��8;|$�pL' ��P�>Q_Ā�0d��a�����`^C	l86�ȗ�^�n��K�����B�O$�f,%]З�p�9���_�z�
�M��Le��>�%WF.^��Eˎ�~5.G�C��M�{�?#�)���W�A~��f�t:r;|����+����$�*,��Z���NT/�ҋ���0<�!>X�U�q30�qKw����;B�ƫ�z4Q�g!� �/�cz���@�/0B#{3KT1���/;�$?�P������37���B��U �"_��F���"Z��,���8��ߢp�w�8+�^a��7�b�g2��w��0����+� ����*��p�Q㓶�,(��.�Hv���-��Ď�E� ���^��ђ���T,�[ԎJ��O�1���=Nd>�'\b��=v���� ݥ2/	\�`��%���j�Ix� Tӳ+8�1�����/���ߨ��M(����O�Pk�jEA0T٣�@盯@Z,y�p�~��L�ohu�S&7���PPu�{��@Հ ٬ݫ-}v�N�d?+�/r)�A�W7��M���,ݭ� Z
�E�LK-	4�+Ȭ_k��i�
��we�4KF����YٜU��z��RjQЭk�,3���9��:м4F��ڗJ��"!��{NK��Oh]�t����vK�2"2<W�q�w��$fP�c&�G�*$�c8�ގ�����ӫlw5�-���� t��g6j����^\��đ�tm��+sKH�W)�R4�2;~����_^V-�A�<�M��d:���m�;>�8`�V��`��	��`� �O����=��ԛ6Kh���h0�R1	ώ���h�G��./���#^&ֻp �=YCU!ry�B�x�ߞ�|��*X�҆-:	v�r*��J��|	z����V�isa�=�j��̴�Y��2=�9�[{ q�ի'��?���)cMl+��X�ݪ���į~��z�j�LAU)1Y�*	M-�BNzK�חWtQ]�A���5H��Xymq�Òy��;�l6��<o��jH��&e���Q�֞�YHu?�'���Z_��Kߌqwo���7*����㱂�W�(���IIİ��j .���>�_
&����MW�&��9i%�#�F؇�Drn΄C�]�U�MVbFqƱ��u"�d��t}���zX��b\�r^�r
��(��$����tk� �Ə�x9�)t�� ��<!�wU�J@���?��f�����T�/�� ڣӚOril}��7	�0IO�;�^��T���z������pnI���o���r���sj񰡖���H	򢢁�r7�E݌+NDn=Uf �uHM��fw4{�~�p��G��&:?�q����*�?��ԳK��J�����`�;MLpy�����9M�/A��b�o��4)��?�)
�ʝhQJ	Z��Cf����:�����Z��_8Q�6�0�4I�M�#��J*�`(	iݱ��kNB������M� �hi8̴�$��^���xoL4�?������8����t!�;��Z$�B��|��z}O��{�G�!͋��:P��tW�a8��Z�,�~YH��W��=�F�+���������U�n(���g ܱ���o��?�h�@��ל�Ay���I~��r�[�{t����W��-��k��d2ϯ��J�H����SF��p���9\��Aj��i&�Z-IV���������ϥ-�|���Aw������ʉ@��F��VpK��;j�hbm����[�	�
���%�8���u#-�+���������J��V�n�j�c��Pdn�/�*�״���X�
�/�l�V��n�%y_2�Qg���11�%������Z��ɨDx#�;мDQC�Zk39��s4�h8�>���2�g���l_�il~=8���23d��$���I��{�H�7�C�[d�Ԗw+�y��V��q��g�OE.�1���O���a�O@f��dy�
hh�J{�8?�|d0��T�@7(�
�Xe�
���My�"�I���d��8΂��[u�?t9�o�,��W�OC#R�6!���˅	�UH�!�l!&7Q8�'�Ĕ(�B빍.(o��&���JH`M9)(�[�#�����(��5�9H6�x�Ae��[T�7���AN��:P���O�m��r<0ՀZ�,.��bu(=k�`T�)ͨQ�ݐO�#������IWhDd�,�Q-���f)�o���Z�^����b�����Z&��q�b"���Ÿs��tn���Y�l�]?��g�S�3-���Kkb�Tz��ɐ)ܬ�ߊYd7e//�BqECˤI�j4z�_Ֆ�w�D�n$���w#ʣC��)S���/�r����ֺ��-Y��QAQ��������}&Op��64(�*��)iz]^Ƙ�sihT���� /DEdwz�ϸ'��"d���֌E�y�<���P�]���ڋ�w,�Ɋ���cZ�6*.!�����*ؕ�I>p�P��6m�.s���/�F�yyـ�'�^
7�"6d�7 m?˚b�7���s"�e����p�;���Pɞ�qM�_�/��	V=�kTHy�&ğ��E�=h�O��F���:-_);���T�Z�p>qbjd��������5J�=��Y���P����O�V�B�mQ1�8��~"�8�N�k����I�+o5	�F�
ŕ�I�Ɠ�Ϲ�{#�2��#��������s?��)qP�I@`.Ұ7S&2�/����蠘U
�G�����.�L�P-��]��[��%�!~c�O�r�9���(+._���6��L��������o��hQ��N��k��7$d�t�ĵ�2�L��~З}L��N��A2_z���@M��]����?󟏑� zx�5��YB~�s�F��L��������Xh#��3�@V����#1��j�](��8p�������q���ss��%���!�����2��+���0G��a�,�l�8���5I���F�c�Ϧ:�YU ���,��~��_T7Ϧ^#�q&�C��ϧ/3����8+Ȳʘ�|�ו%e�I�e�7�4�l2�(S�5I���2�켧!v5�0���磮��u�ӊ���p ��vq�hb������S�y@�pi!~�(�Ej��K����$�x2���
�6���8n]GL�͆��ق	��<`�T�8���C��w�9]�B/M� ��m0��e[U�������(�|���8 �3$Bo �����R}�+0OGO�Y!���W(b�%W$�%����R�j�$5Fy�˦��s~�<�21��`�@�%��[���3�b���ʪ�8_�YY��]���㘾�46��#Ͱ��Cu�e3{�v&��f�t��t�|��dIǫ;�d��7���e�颸l>ipw���>&˧�~$���~@�7���x���Y���/���U��5cIv��/�Ҵ�5Խ�$Cx4�� 5N>�#���Ǫ Haj�r���6i��s�b���dC�
M݊�-�Eq0�K��o��q���T6���]o\�%^KёN�A��d�_P/��X�g�
@kQ$����2�8���t�k%JF6gЫ����v�{)��d2/�R��edT���ثx9W���ѣT��~����'�D��-+����b�b�U�q�Yu�p[	�g`�+f�v1�ie�9צ�����$��ވ�y�3���t"�gO�t�VS���x-�z����|�����вT�k)��6�!���ڣ@#��\B�-�� Lr�(��#{�����O�l}i���ܳ�4n�ފ�I%^�(��%ﮚ����Mi4�ʸ���@���sɜ�nZh�K���� �0�6����_�	>�ۧ,�<�믯��(�g�̮�?���V�|jd��6*c"��� �w�&��A,i/�r��}D�[� F8��8gKQ��9��x 0�:�=Jp7��/8��%���v2�[��Q�f�t����(�Q�$�\@��*������~ד�>�Z�22�T0v�,��5�/N�Z��+�G���a*� �ӗ=i���`�q��z'��R��.�7���l�=�3����f��}���G���hDt	�ob/Ye�xI���oq8��]:�a�H����Џ�����/�cULpv�.�c��{y�'ˢSk���Xk�%R�]�9�k�
t�; 4ek|�x:xh���Զ�k���;PgW��OS!V�6Q�?���� ��s�A5"U����ߌ�Y��2q�ҳɩ~귑Q�6�[�>^�h�L*�T�pG=�v�5�	wU���SZ�HE�W�y���C1f]R��v��Y�0��5��| ��|�B���z�F�d(j߽�?��k}y̝�7�Ȗa�)����窪���h��q�i��0��(�M��mMtA )�X؀=q��0`ϻx,3�V����-Je��L�;�8|#Bp=�S���f��''���P;��ܙ����u+�N����	��OOhc��,]'�V��<��ײC8\�R����$�R֫Lͼ��؎U�a�������y:{կ0���Qj�����@o8 ��0�ɸ�N���A+�I/?A?��L�+	2p�R$�*tj
�2��ud�l�*�ZumN��(`I8T\9 Tx�\���_8�7��&�h���
FRl�ŉu�In����O�!�r ����7����<�_�wL�n��ڏFK��,R���ҋ��+Z
Jy(�y��po+�y��WWy0(9�÷���O~�dy�%��ʘ����J��:�2�`j�;z���#���ig
�lM$'d(��X\q��8p:s)Mi�f�&ݵ�in�`E������}J���֯�_�Y(���ܺ�Dע���	Z�f�}r.���y��V�Г�d2�yi�O:�W�o;�2�t'���rJ����� >�������䷂�����|Io���,=:u����*���� H�RD�@�e9���!<�/+�?�R�GhZ�%���Y���3����s��{Ǌk��k�M0��I��%�֞T�c/�YL#�u����5��hD�-�2��(p妝BK��8�۴�yKr�и�R�	>H�jp	c�0�������M����Ո0`7G~�^��m|���0��|S��an$�I��Q}�m�X5��H��V�ֺ�b�l��o=����*�p�uݱGT{�V���.P��o8��Q7F��g>����T�ΘWjb�9��R)��;Ws�đzmSG����D�k���G˸��:s�Ӕb�(��N�����ں�|���D3���k�P�!�G~���� ^�W�g�kDb]'A�)�����,?T|(&˷��J�c��46�ʢ�vʈl�Q�� 3K-�մ���T��l.w���#߆�@��#������v���w_���h��UB�	<�jx��<ڜ[cߤ��I�Z�����P�l��1�D�3�<�2ùP{�ј��'M e��O�:LMP�hJP���T�����d\�h�w��7�w����'�{*��R �x���V��豪��<zk8�E�2K���I���j�_���R��]����R�������Aҵ��T�<�ޯe��%P[�5-8ty�ƢE1�B<�n�߹fk���\�/���[�@1a����]Y	�)�x"�Q"wW�(�R��q@S1��]�V^���qQ�bSW�.�(_���L;8fU+o��H�-"tr38��\��a��)���~��2�ƶ��㧞��P�5��	S�u\�kyr��qb�Et��Cr��0}O6�-�^�x�ӟ�3b�#�� UHUQ��D��WJ%�
�۸������u����Y��X�'�`���br4�rG$�O��g6���S$#��!�0��Dō�ք�#�4����c'���GyW�|��tԞ$�+{��R'�y��շ��m�مjD�u8Gq!�����x�he�Cn��`g`Tڧ�!���QU�]?dJ�ނt�����>��"`B�������Z�
��V>�^
����g��f��ң���g�v��v$�4�u��3���U�r>y��@��I](�)���<���lz�N��|�TN� l�{^��,����V�ؐ�9i0{>^�a� ����t"�.��:nbSAj���lX��2�`�!�-��F���4`�������[��b�ވ�͂�7+�ܬ��)�j��-<�ԅ"�uZ����R��@�*��4��,C&z�g�3�C�aB��h���=��K�ٷ�A3eZY�y�67�-����gX��p��ѿH3],����&�:=�c�����"�֛�< �ܖ�ק�,_G��2Ǎ!�-���Bq,R�N0���Bf{	XLLy��1�@�
��uɕ�F	��^��n|7�;&�����2��F����>)�+E<�@�t�8B����er�(q�4��UG��ߟy���R��]&����Y�X�)�Z�~8h	z.��;�-���� SQ�l���,�E��m3��s�O��rcGJvq����ت��/)����Ӧؗv�,�OU��J��$u.n����֤����<�y鼢�q��My7�I5p�&��F��n�Īt�<�N�<l��dfgI�Zt�Yz~��k"g6^C�=�4�Hɸ�I�T$X�G�������~eYg�H�m��e@_�!�Sf�����]�ͺ��>�� Q�.�PdNs��+>����*��&�-�ZuĒ�X��B��"!<�19@H� �"��i�ɧX���u��v�%�ߍò�Ub,��A�������]$�+�障	%Z�û�!A�}�т1ͽ��#�o��̄�*�	\vKy��w�1�35����ĿͶ�u���#$�f���u���Y�@�i%p-|@V_�šY��c]��l����5;���!CD��i.茪l/�6s���ů��y�.��A6nJ��w�vl�pU����Xv6���_L�̫�����/J� 	�gd�<,��[�cA�����aM^(�	���m�G�cyX�t$�vd�_423��I��&�0�xn혿�⡶H�|��m?��#�
�����S��D�5V,'�q�w�*H}(0�JJ89ۼY^�vr��.��~�ýӲ��{�%b'���˯��aG����]��=��K�A<�v��S��V� ^Eb���#��0��`Md���Y�*t(2�̽n�������βi{|t��"SB����YCIf1�=��8�K�!���D�D�}AHV/(KY�#:��j�_\�.��EL�tĤO�ṕ܇�"p�s�+S�C�Y�*z�c�^���!���}d�������%���d�snH���{�� q�A2u�;KR�PH�#V���9�"�d�u�8���?�Ыu�>��y��&����[��0: |����h5����J���˿_��Þ%�㊈��
Z�Q��j��q�W��ܰ�_u����W��p[���DR�_>C4r��`��HEg&`���e�C��\(�I���H�=j�Y�W�Ġ�UC�'ԷV;�'~uWqz�Az�\ٞ�=6���8]C�̓)�'����9�,�5r
y���:��3m �%w�*�w6�/�e*ȴ"9>J�S4�/��WjU
EaЖ �0����`�"H�GoK��5w��fb���`gM��XT7=菟%49��@��o;��Ot^YN-��h	�">y�v��z��r���$Izf�dd�^Nv=mEKځ(@l9787@`��D��j�z5���Q8�&�f�
��I����Q�ڛh���0��L쐳�jp�>b�";7�����kep�P���N��lQ�ݳ")�(Ql��)W<͠�SP�S�m&
�[�޶�\���n�>�=��fD��.���4�5lJ0�^K�$��X�"A�c�G{T��>�2~��5@�w�SE���T�)M��O�~����v�/��)ߤ��9�A=��k�EOd3�WVT��执� ���|��
M��-�F �%����A�Aia�p�	>m*���I:[��;95n1-���B�v��1�f��}� ��(z^$��m��&(�P�U�X>�I��dudo|ߦH��5��~=�Ы�)"ʁ���;�޲��U��OTغf(�i�)��T�w^������L��Q#����v��	E�6�z�=?e��)�ڊb��������:{r܌��z�D��\x�E��Q����J���^G�T�ѓ�̞���t��10:����U�v�?��EY���of��h�y*�]�Fe�˙�2O���h1C	��,l�=G�r�;#���_b��RC9������O`t�N��-5���eD���C��.�v�L<x�+#��c��?���Q0R�u^O�Uw��	x1*�ʡ�YP��I�R���Uw �j��l��o���5�U�L8�쬿M�Ol�O=��mH4����t��Y�ݶ|��oN�u01�i.���}���G�a�y8G�>ѝS���l\3���6�'	�F��O�g�vr����q����<�&��l&z��#�߻��`��K��}��b	���I~�¡���'��="�T�R4��9^�u�	{pig����vw<����r�ĩ���i��,+EA#���!uꢦ�������cKӱܭ�X����4Fk���������!�y�yiw�	Ǳ�J@l�ܖ��d1�����-X�D��m�b�7앳ܸ:V�^7;� ���a�2�,��t�쾉@m���Ӭo7��L���'�m��qp&�ht`����}��S��2�Tp��/mb���$���x�9��� t��;)@49��
P����ʫ=k�[���r�.�T��p� 2�;�hɩ�v��s0����.���(�fZ|d��u&��j�\|���kS ���"OÞW�#��6t�"�뜤P�+֍ԎcQ<��%&��A
�>�{�F�C��]�:�N���'�Q#I���{��)-)Ml�G�XOPpyY���Ⱦ���*���:1P\U����80"����qb��*�����.� ����2��\�ʡTC���?WM5�g��J&��@_f~���Y�mG�%y�~�m���ļ;Q�>�גv���hև�d�\92`��kU��U�t��i���x nJ�q�4u�o�a���H�[⭽�sp����6*�����g:�b���� �o�k�K���c�T]�nl�aT胻��X@���w�_��H"��~@�^��Ȟ�����S���ұ���#ҕvp`�ի6L^���h��²g$����2�Ւ|?υ�@���	a�*��"���W�+<�<�z��֫��wrSW�Gb�ԈZ!��Q�E��ڽ&��p� �ΐ���NW����m�I&p���w�ڹ=��RL���Ud�Nf@&G���d!sS�Z��M0(�e�$�	"�&�=G��B� q)�������TF�����4�"O<ţ�.�6�݊���Y�����0O�I�Oc���m�}����≞f��p�6����xhƙa��|�+���Kc)҂�Z���w}���]�`V�����W��a|k��v�7���>5�c�1٩8m:����#3���>�5HEs��ՠ¼:���HfޒB���{��.vI{~!�i����B�t%Q�`�!��F�f���������/�rj���ʵ�4�1��?�꠆��F4i�?��M�Z��ک%�9ء��`P訐;6F��R�w�P�,G�Q(�S�ћ�\����ܔ�����K!�F'_��D�.)��W0���͌?�����e6�_��eY�Z��86
����NWz�Y��,��
?�Q�I�Y�IM��EB?�2��Թ��ε���5��'(�>�_0�WN2�:=�W��@����oN�5[��g�fۢ?�e��K�~-~�%��.��H�}��z��^�>��iC掕,
�ʟ���uF�v�oOs$������ ӒHQSd��dغ�Ew�9�yJ8Ϣg׬u���6N�=YX���̖~(�x�Lv��5Ba�)��!��m��*�v�o]�d�F��:C�:Jxc&���6��%�o�WoQ�HH;�����01-ǲ�q�?Cx���f}ҬV&������Qui�1�m �Į�y������Rc��Z���YJ�-�{��:����i�y�]?QR؝���㖐���.�R��ͦ�<[��j[ns&���1�3�SBL�1N�'�h��W�x3�{O>��Z�.i���kdʢ�`�rФ�w�j��
�1_Ì;g
��Q>�qR�&�ɠE��|pw�ݤ ���,���wl�\k��@�в��Ձ�ckh������g��r�����[^?�-D�ģ�w�>�[��H;��O����^9p?Z��YA|��N|_v�/;Z���2Z}�2nJ�~O3J&]YI�E�O��H���.��\�C>�cP*^������լ!z?k=C.��T�#
��-:�r��Bo`	2��}�����?����Zp���Q>ˏ��'vDe{��j�pr86)����G�#�ķ�;;jƨ��A�UѲC���	��*�[����d��&w�%w�@�E4��p�� �$�t�������/����R3��	lQ�ޝ
F��J�� T�
OE����s�����6?�j�j+�}�,��_��%d�bB7T&fxI��pՑ�#��r�D@��C����b'��3-��L'Iu2��|�*F��`�1�U��2�q������ŕ�(�Sg��thr����F����*���.���%��:�準�Z��eO<��̚��!V�u���k^�q�D�,���XK����Pb��"U�#l��B
���;V�����Rs�<�g�i!b��5��N�{9'�����
r������*O#���4}�Q��R8tgGj"4�~�����{�z�A2�sk�A����j����pa^�<����HGOYA����]���U~oC�	}⮢� H�s�d� ���-�gGerp�z>C3*��iU�=��*�i"��YYEL�D����;�pSs%����� �'e�hئ�y��Q!;�G�"OzHZ����s�Yߟ��Q���b�5� ���6�j�����bW ~��ǳ��m�[I$��e��6�P��I7�G����PΩ�5�Q�����;����('ٮ���ꐦW����+3R�g4��_�\>8�v����3'>�\r�T��Cѥ\�����x,@Cx�Z�}���'����M�z!�v~�Yդ ���7��p�&JV��.U>���~8��S|rg�ަl��b�T���4	.�ьm�(th�����Jڼ�dD�_�eW���o�xDib\!���HQ�!XvlH&W���:\���"O��B.Qi&��G��Эن��W�m��P2�[nx�����#i^�3�(�)���ثi�x��C����;�,����v�Uy��	pq��2���R��&�-30f(� ^���K:����p���]"Ӝ^
6ZS�)�M����ׅy6�_'�����_0D˲pe��_?��Y�<��ۘ�nϸ=F1{-���ip;�B�8W���p�����Ц������ꖝ����w�< `>t/r���6Ĵ��@�x���\��;������*"r`�h/�A�Qd�q*`�G�y�����'�řh?;�Y�#4�zW�	���9�[sZa
lac�jK�&@��+�<v=���C�؉@�7���+0?�����yOR��%9�I� ��6l#�7��{����N�)t�B�G�&Or4�>=�j`�Nq:�@}#�h�"(����`�_���5����n�KQ�I�>�T���.rkי����gN�ޚꝿC����ٵ�!Z�&9h��Ջ��43r�t:HU?�X������X)QX��4���l��W�+&��UzDߢ���`�B?]�ci_�J��%��]y�H���T:�4j)�y�=oE� �1"��2��;D���Xh�&os��,�`�H�Ds�w�t=ۆ�un��h�ҡ������H��|/h��F✔����QL�n�=�*�M������Ut�zՋ�C�����j��VGx�!$�шA!���,nGg	�/�^=��EȆ r��rE�)�@ j�Ff:�lS��(�#�,M�9}���s��b��;OmJh��3����^�
��b�if\��l�X���A��Ud���n0���s����o����	��-Ub%��A�\�UB�7E?4�ْ��=f������7�N���
,���B��&��<�yu�<oo�V��A�o~gtF���TGZ}n�]���E��v���)שּׂr3�#G%����U9^�a���,d=3�Ay�
���n�?�r��RN��~��X�S����uYh�}��A����>:��H��^�s=6���d�0k!'��I���Q�������a����Zd��x4o�ө������R�iq������ή�w3�hL��b��?=���w�T�I7��8���Ί��	6<U"ʮ�&$s;��A��d�U�6�F��٬J���%R����Ͱ5�Ӹ��CA>sW�����W6��V�4z:t|�>����]ϑ��n����?/�	!ֶ�R���=�"��4qڐd�dr_�[M�1�C?����uF�*����_P\���AO؊T]1�S�'X%�(��������4,�.��h�N���|�ѳɨ:��c�5א+Qe��oP�7%��fg�'U��a?3��3r7!����)h蛒<���E���I���J���`	O?7Hpid1�+�EΖ9�3�����Fr�p�b(�b���[0/����84uϯ+n��f/yN=����!G�1P��r�XG�C�_a�դ�sո�;J|@~�e�BWq�?�aM�DR������>7�����zV�(����yJ{��V�RaF7����.ZR�@���nr�d>A�\����ؿO�X��2�a_�_����8�=���#����T���񒞮ʃS��I�T�N�"ľ�������pQ��]t��'�YB�an��Bv��o�����r�=��d�L�Z{*�n��E(����g��W��kh��J�%	.�a��G��[E�;��'w��O6zW"��.���3`��CP��#���n�7�Eg�J��Qȵ=�|���pְ���g��O�>r���$ǎ�ԯ�"S�����8uRL�$@��B��y��Jj����%w�L�����Z����]�e
z��b�Vv��_QOER}fX�D�:���>�IHO9oP/����;S��|��u/^�9�쇷����bu�����l��l'��]��`tzTV.zU+'�R���C�`��(��n�V{�s ��Dtg����ً�ߠ�k^+#t!�/�p�d�)1]������')I���	�2PL�5��
�&6�6�;�1��3HKh�l�\����/ܳ<b����8f95"=��Y����?\��4��by��lCAn�f�>�ӿ����}���+�or|K����ZV�@�!dAw����ǎ�����>���H{"0���Yᵔ�ֵ��_����
�7Rq����.V݉Ax^֧�}sғX>F~��~Dz������ߦ���m�;:y$��p�t����3�]����d�I��9�nI��Z���"�V;��f
[����v�ц����TE��Ɯc�J�75 ݩ�ɒ��9�@�tt�ق#�D�F��胔ٝ;9�ЈSqtzmKУfT�� �㔟%rR�VX�Z�C=��<rx{�9��s])�p)�z5p�	VUJ��pu�m�VCfU�a�F�3���-����%2C���K}ݢ�=��mY��2��-N�w��N�"�J���пe�,y�y���?������/lFi�fLL#�?�kd�YQ�ٮ��ӣ�[���o5(�	���3b$R��X�{�M�b�n�q�\��ol��f�6�*@,5�mh���Sc��nH��#w���Ruqv�,���pwRs�Y�/.|b����l��O=cܑU���@]�ƴ�Y�8u�F��-��d,�<㒔t��P��.��8H?�!Ƃafi���Ag��!�
]�7���%�!pM:��(g٩3�K�T�C�.㻔 rA�w^ά��*0��-��V:�[D���0���6�9��-��qc~��?���W����r6KX��q�����j-j�ο���Sj�Cn�L��(8������#qƍB�ՏvD�`X����#ד2˾H�J��C^����m��z�N১�$N �Zޙ#fve��O��[Y~�>��o��О��-����N�[uv	Am�Y��lB�w�3v�����ݪ�a'��$@���ߛ����))�$�ad�;Ì!�$S�p_<-�ܜ�k��euc�>�@]FTV��Jd,�XZ�u��%|������ �	5m�y)��u����~�=x_o�����32@�,���]�|���������Aؠ�E�r��{iv�x�w�ȶ�^a���h�V�X>��⫹�dp�VA�D-^b~��,j/�m{Z��X�ֲ]V�w�����,�L$�l�\�B���4=�Eo�⨝��ʚ�'70�9(���O�	��"����]RZP��ѥJ�>��Q6(ǋ�73�/߿�Sx\��B����8��n;��{0��晦+4���-��칀��=�f�Oo�?X3�UF={�2N�C�!0)(�U���43�X��Z��"�TI.�� ~��qz�{�OSY��m�UȨ���d>j(��<��WT��\Ѵ�/��!����Y��4�Z�\y�
��d1>��P]�^j	�Ʒ�zԁk�\�!}YD�EC�9�P�=lA���A\?����6�Sj����쿋���2������D.��1̭���{d��}�c�2���Oq�m��T*V�����O�1%O']E9���0�>M���l;�����a�c-��l�&�!T?С�
A2�:C�d��kc�v�︪�pب= c ��;(IM6����q����gXuWr6�w(,���b|�B$k �Tʩ�%����d�/V���m*�W,��w=Uh�
���ӭ�Q�����G�k�Z���7�汿֩4�S��P��������w�KX+�x�8L� e�-/QW��6���0E-��Ui���Z����Y{J̣@�E9nP �'��������~^2��:x`�}�ʽ�抙n������ac��}�Y���ȓ���Q��@�x�t��z{H�n�L�6���I~�Eu;:3c�]c{q]�b������Vg����m���U���u)'Is�vR�S�>M��ى�~tq�J���'�q�b�Q��aޢ��d��z��Ł��}lH;��a�`_7�޻�)��}d�\r���62U��>'?�Ŵ�TS��!qf��]���o��5@�z/�fa#�=��l�BkL�Y(,dI}����´�0���edg�t���Kxe�5,@Ӗ��:��5��QH����D���;wtr���Z�)�*�̎V�
���0��eA�@@���f�2�7�h�a��\Wa����K�Z�h��ҩ�?y��a�~��N&%��9�L�[���/s��v����������AW��a��j?d]ӑ�!���k�����@�Q-�{�l���~�S��mr�h����������G �uk�Yt>S�?��n��H��]c�dX�n�[�"r�iJ�]��I�"H�|�Tl�޻q�ex1��xW�L8S��k���/�:��)��<�*��&S�! ��Q��v���Д�&}�5s4����Xݟ�)�,ʹ�P9��3�-@4�O]��#���}��9�C���ś��D�j�W6��o8�M����O�tB�c��;dt��a9g?�+���G�3 ��;Bj��&,to�:h��?��Pr��I 8�!�<�s
��⿿��7�J�	�g%��<r��	̜�M�+����2��=_[�Ѱ����D.�<X3(�t��fg��>�I� �#��� 1G8��4b��wGK�D���j��W�)���}�?�UF[���J%=���̲�a�o�U7�~$Nb�Kt���3/m[bS���rc�~�=՘`�t��[@]�}Y z�{>�iJ+_+�R&$����j~�%չKC �}��q��M��TF��o�O���7n���R&��g���MZN��ߍH
��&���T+YE��?�퇯�A�ߙ��H�t�����9��<L�"0&�%M�2V����e���2�c���h��bВM�C�V�ˣ:��͈�6����=)��|�;�O]4�R�'V6�
'P�\��]�P��j�a���U��jC����$kb7��z�
�{-�@Z�QisK\c�f�
�!��#'����l��9�%S�J�(�������t��L��,s��z�~H���O�gp�R)��ө5����pm���Z�WYɫ�ܵ�:c�M�AW�\��O�;�o?�?0�3��<�4B��<�J��W�T':�<�-��P�9P���߾�&C�5��������mZ������1��T�����VMk3����!���9e���0&8�	 0����6�Ƭp�Q�*��J�8{+�&�i\P�ϳ�!�&�n��#� �y�г���`��7S��7bd�֙W[�%Q/*���U���>����k`n��12�TL7�����n����J�.���,|�VGK
����"�+�*�|B���/M�hY7�`b�S�u��5#����nLi��C�Ϲ��L$�H`�W^�"6M���
Q�����F�Z�duF[�)���L��Fc^����Xx �<�M��^yEil~��:cl����K�:���H	{r/|Nԛ��3>8l�E�<��-��DL=����G��J,�ι��.1��������m�c���Q�	�e5;D��j<�.Ҫ�t��YTĕN�����3�G����R)a�0۳C}�bLY�:ND��j���TC��'�@�����ĀI�p�9F�^�twJ���=�<��898̟y"K�����_�����p�Q�I��LE�3�hr�<"b�J������x�$x�kcÇt/��5�:a{R!��Y&�~{|� @.�qLl\ڰ��BdXV�K��:zyJHIVZ{���I!+���5����o���*y�v��~Vfw9���e�� ��T�MV�Q���t�^��C����A:��A�"���S�iV�&�L"X�����t���?���E_bf�&7:��C�{bEg4�;)�0��%Ǿk��5���U���]س���q�hi�`M���iY�ON7X�<hW����R��Z�_�Pn�P��V��H3�������T��zL��h�9ri�<�('k��Z��f<L�i����:�a
?1F>�ǡ�%���)��S�w��0���1;� }��D�:��t�V59^_������f���:�W��?���.*݁5�eEa�d�g��=@�k��p��Y�"��{s��@KǛ��9�_\J=��Cw�����M��O�� ��7�iy�4WYIl��> |Jy7��s����"��E�����67�t�pcB���qX����p�C�& M�e�J��Ǒ�{5}~�ҟ�U<�:��Rr��=Fe�����2,F�����z�ƒ�uT d^�&�#v�fU'��WXk�5��.��&7�TR��EQԗ�_�2���U�B�Y�9�n�T?�"n1��/�L8��*C�j�-��V��������>��o4���B��<:�5k��,��x�%La1Rn#����\1�^>��
��̉�*�D��KթS�ʮ,� �gxk�)+|�?��[��x���ԛ�x��o���:�{�Rt�P�$O 	��Ԡ��u��Xӛ��������5�ع����=�}% <�{jd�I<Y���������S����dN��fa!t�6���\��:���H |/]6�ad,��C�9�t���ƪ9�o�nۙQ22�=��y�BaC��U>πa�$�݅8�`��������Y�FZ�{�&Q��a��x#nA
���dG�$��U�|�7}��
�� �ԭ!�����3Y;~�!�E	MպcRD̟�<X-c�<��G `h�tƺg�L3M���-�T�a\��x����ĳIÌ'��`�}��Kuz�����&"�P��Gc9cVM�O�������܇�R�ا ��Y�b�����?T+�q1��D���f�\/A�h�O� ~���e�
��>�V)��&��R�qH��R��A�D;���OA�>E"���J^'��ƶQ�'�`ə&��
&�lt�������������w�Q8O�;���4GeX�j��O�oݜd�北�k4�ΡTyGˑi�vN�F����fp�7d���,��i��7����^r�£pRnZ<	��Ɵw�^A*�����a�N#�w�����òI�Sm�9�8͏M����W]�K�9M o��n��oǝ�]�c"L*��f*[��t���{8��-������Q J�3�OrXy�v����s�5���v��U��j5��Քp[�ј����`D`���@��\�E�W�J��(����y�ΉPE+\�8X����F�?�ِߞ>cV�v�do�س�{�O�%5�۟� �+.'�*�Z��+_�ŧ��3W��Gz,�: ��)�r�8�'�Vq�$�V٫O�9��~@&���řy<��m86���{ۭ����hZ�`�
��I���3=� ����{A�F����ɏ��r��
ӏ��<�˞��f,�y^~�X��w��S�T�h8��PX�2I�i7���nY��-�����7D��LJ�2�|h�tbl_ob����"���R�(WcEÝf��_6q��",�Pq ��������d���Ĥt��@/{k�(8B�`�پw���=FCL�UM�JL� ���"ֱw�6oW��ℼ��O�mP{����W�k�k	�fh<���=�4x���y�Ch���C͇��&4i��ü�fg��O4�
,����Y��\�&̾���l������=��ֽ� &����D�,IP���/�nܕ�+'�*�N��F��`o�-;W���b�#^�'}���悒��q���o���\^h������*���7~!A�H滑0�W6IB�\7�Qr����i�I��T��of����,F`�.�WR_�8�g��,Ϡ����ף���#��
f|��+�o4�k~I�g��`�/�sj�_G�u���;��Ig���1ޙot6��D�X9�4�!��E�a1�ԡ��z�?��ug���sN`i�=�5ި�1#O΍ �E@1r7WVVQ�ӻ0u�����Ƿ���8�L����s�]�o��k\�~$�[J��lTj�.z���-Ҳ��'���&�RW�Vn�}�I���h��3\\|�9�p���-��`�M4���t�P7�X��!��_�4�l��_x����-!=s2�7���|d#a���>�����2����9���gƿ�XQ,�b�.��Sp�噧�T���:��d�ԉ#�D�`��6���zB'e�&�i h��r6��k���>�	ֻ�c�Ro�%ԪɅ���hy:Y9��3��N�$`S�ho�$P�d�$���驁R�|I+���S�7z�X�z�ڷ0�D�@��`R�Y�&��VvJ�י�5��$P�����`��y��kI!0���F�̯�/���E%z(Rp�}˘gK�i!�мl�n#~��0\rE��-��b�~T'����Y��h�֡+��g� ",x�C���x-@�'�պ�q�2n�tZ�X��0氫c���)��-�E���!�X���/Y��������S<��\*�N�!���݃�� ��If�"���C�9����D*�0(��**�4�ucO>Y���Fq&�vL���"��P_�j6���5)Z_\�����U�L��Q�c_��g@;���K�?�C�e_�la��Q�ىSN�7X��M��^��bO����9��.3��"%f�@���a���W�gS���s?��,�V����}h�D��>����xU�XO	GA�#��qI^�]qw�UlLo�PD��R@�����C���7j���h��=��alB.\V�Z~�G�ys��y�b2yu"�po#�
�7����������� �z�r,��`!輝��e4V#Xzs��&��֏ 	)$=�ú�a\!/�\���uưc?��)����.o��l��W�h=���!�5萵r
�9��ѥ��o�TF�}.�r�L����z�������D���Jr��1��1�������}±����ۇ��g���CQCק�@~Y�/�6r�8B'��',�v^�\U}h ��J0FK��Y��*<�|_�o���*
=�G}4� Қ�~B�<���E[�8��1,��F�G��9z�m*�+P&l��"�D?������0�;��i�3L���xr���!7����'Qi,��?�����_�>�n���$�'��&��R�ߜ�$�(�k����O�>�o�{w;H�������U(n�$��Un�$z������D�U�]�x�Xt�l�U�Ԙq���oW5�~���s5�n��^߄;�@N��R�+*��{�ݒ�n
\3'#�D68i�aXw2]��ou�>�����t�?uT�k.�;���y�Zk7j"����fI�c���-�d���kl��(/���W��Ö'�d��+r�ss��P���N߰�A�5�MG�V|���u/)ZHvs�ZL)�)���~N\��/3���G_ߴ���Ǹ�f#�پ�[[���c�L�Y4�ۣ~�T�	�zO#��� Ԕ>W���Ok����q��dkF�W-��"�7��u���SҞ�^gfߥ�gq��^C.����������Îc_y]H�[vW�־��b.X�h���S������D�V��7<o4�S�����Y��L����;�)rZ��ϒ�U��K�{ȼ�o���۟�*)��	;��k��O`����$�l4��+q��<_!�Lm2=�L�j���.?8>ù�U�3x+�k-�?�9%�"?W�en�e	+ �9\~����]C$�=����ж���E 4�+��(��p�JrL������
������gW;Y�"z��t ��O��¼H�$�S���$�8C��8ϑ�cs�=�C2�ڭ"Jo|,�����Y>��ֿ��A�ltK��z��	h[x����;O�	n~��PA�����"�f|��s��N�9Rɣ�9���Q�Nջg7��,fh�U}���b��bOH,�
]�L�/wI�Y����x��>�zx]�|�S��  ^�خ�u���ը�6�"c�	�_���#����B�^b���q��:&-]�#bXf��=�6'*#�M5g%?@&�I������I��8Rp닲f��n2�I<�=}�@R2{�"��Mҍ��p�#�@m���ER&��# ��12���IEIf�YAl�D�ݍe&�R�NU9��}e��5=������HZk@�/����4W����-̓�˯���|g��Ew����{���q5�U]!�y��g���ccT�)�Ro��v�)��,BA3��XaO�%8d�9N�N�u	j}�ǭ?�����S�(~s�(�L�M������^"y�^p J�-��2��/ɬ�J�SN&��n��6/V7s-��,&�o(k h$��5y�w��^�tX1�G���Z�˹���l
��W�ӯ��`���o�5�)��������K;��&5s@O6<HyCMK��s<�m��ſV��-ks�����fn��C�9��R�/@�������L���b'�KʑZ�;C�N�F�P4|��X��#�X�Wr��i���}�.k��X9�[mz�U��?�C��xl��#�]�:��H�ͳ���8�YN8ڢؽ�4�
]�M[*�Td$�j�����6�@��]�gj�7�:�n�T���#�>��*�&n�@�S�!d���������%�(�]�
�	��d�q��1K���	���]�m�Q�ZC}���9�)�=�~%� Ru�yhLI�她�@E��@n��ml�v��p7]KL#&��ʭ��劲y��k|I��/�>D�"��^SB�@��U8ȑNF/%��-�;�o���4���߃�hT����8�%'�V�>�~�Z�r�����L�gK\�4�e�P��#�������TН��?����6�&+Sz*{zx���lE�񤹠
�g�v�&���pOF�AR�
��%�r�j��:�_ 0&�����wK:�$7@� �h�1ǝ]k���8�%r3g��y:���k~�	v�o !C�^�4�|sqW�掝�D��޶�O�~3�\��6�D�ƣ{��oЮ���f$���#�J�sO=w"�̀7�^J�,'�F�=|�b��Eϯ�Ȋ��Pu��5��H2���3��H��V����L��s��2p'	Emd�[�|�fy�zb���|��{y�9t��,�"I����A0V	�5�*�Q���a�l_��vT0iӫ�9��{4,~����_�"������@`��������`"����D%6�u�p����V(�Ν��=Ձ5b�I��6i���iI$l���@&�MZ���˹�@G*�>��u, z��G��"&�55`O�Z���[R%T*��迼�1�~, ��FdIUڪS[��j��Tſ���^�_e�������� �0�%?G� �+e�q4�	�-~˰����i��7uQ�l�:�q��J���̝�Ӗ1�������+�In?��4}+W��q��Q��	wq�o7B��
��+,iv���)���!53��Y߱/���!?�R����_���oʷ�x	���G[w��}�^;vF?��w�c;T�<ؿ-q5S���`�x�r�Uk�x'I��-;X�u���\J"����$�E�>s9|��S\�7�%�� ��|�{��𒉦}�3���@Y;�Jr�uF�A�?f�kD��f��{��jS�@�s�Og����x�'>���PD�pV��H�#�P�*䘏J��H1�/�;(��؟�WJ����U���~����3�"��8`PTz�w��~8ԐC��7�۰��XS�"����T�E��H�åN��S@�ڋ!����#��"(~n��5�=Ek���A� ����X�i �+/&�;�]Ѳ�).��0��j�8SF��!}1���ZD�&bl8�B5T�E4������(��Ԙ��r�C�R�/�[A���)���^D��8Kݶ^Wᵙ�7����x�d��rX�/�h��=}����~H/E�8�!~�<,-���K�������4���(�)vx�.����՟+��5�B���r����E�j⒞�?������#���f9�ֶ��ĵ������@� CMjQ���8���Yٳ40�9a{�l:^�Y
��ђ��L�4�>&��D9W�I�d,C�훚Ϗ�GC'+���ؔM �u\���S���LR�Mo<r��?Hl|>���f�ǔ6�4�=�J��)>ȁ o'�/�0�C[� �l�#�X&��TZ&7�?ǀڑT�B�:.5�����=�$�zn'I&����3Cc/E�4��r�0���7a���y>Qf���g+5S���:�����Iʂ���|@���,�^4�x*xt[Dϙ�C7�L��z�?OR��)}��@NI�-�5;�`�<�[�2��.��i7U��C��k6o#"C�C�G#�|1���@G�q<#X�5�l���l��)x��<OF����A2�3�в\y�B�;�<
6Ng��D�ޭ��~9��@�\�;�Y�X���U�"J�nmV4�,n��
���P6�[���2���@�T��4ᕶv�W\��/<�Mgҙ���mv[�3�>k=�V<!���Vw�ed �����r<0���zzr��%I��F�,���غ�a�n�M�w�o��F�T��vk���a"5��8 �5U�Sv�s�F��$/W�p�f��**�T4g��
�#���輪�6R��+����f=��^�4�4t��Z`��E>����KN�<
��E�b�>ݬ'�n�[*�g+~p��=��0eX<�쟤w���KJ�D8�F��t����g$�T�`;��8w�e�K�ޥN��@��%A�H7\F3���Ae �� �U� �ڣ��0E?��Ǹ�I�;%[�6V�*1���Ò�.��i�n4W�'�����2`=� E�'K �Γu�yJi�m�ո�H���� X��;4��{ ���8>/�K�}Z�.�꒴
��̋�E��~�t���	�q�h	��!��-zf�?@�:=�?����B�yb\�����&U�(/���Z�Hn)eN�z�k�#=�ك��"��H�V��bC8u��������܍�����AV�ys R��7�Tp��%�hJi�棔����<��o1�$t�T�x�Q�Đ��g&��n��}�ٯYۤ��>N��x���1W2�~L�M�����!w�^}b�6�'|��J���Df���8U?B[څ�dn����)���?l���*7�(t��-�)�K��1n�~J&Y;ϸ���6ˇe�9�]��w����<B_�#��]}�һOu�{BP��:�:� ?���-pr��wG��E��UnB��ܳ9�҂���AT����|��
��1�z��T��]�h�g���P�]�1^5&�µ����1�T�j��ǖ(G�e���)}j�T��o������nf�te��v(�M �(V��EϱA;�:��B6�	6~)/	�1�,��Z���s\�W`��c]EH���33���E���Z8W
u#��r�53Sx	LT^�<EUAf�U�^��'���d����-XN����n��d�Ë3f2J��J��Yo�ɾF�AO�����[�;-��}/k���$��+�V��*��Uc����HKY��7��[�Xj�Gv�KP.�b���",�T3�`=�F}�҅�ڂ�}�$���LDwK�/X4/�.z1���� �{C��^>�4�m}H�G���"���%A�M�P��&w:��� ����˭Q���i"a�9[�*:��s���p�Mio>�R�Qn]��6��w;�fap����ji� P~E�	=���'#B�IʀD]p(����3-)K��J*@.�qh��:q�1��(���0�Q�t`�X�	�S��E-��S���X��
�|�Ls�{�c��# �o�⹽�0�
w~�P9p~�"y�+�!��-\l�yy�H��Xe݁�Xp[)�ng ���Q��F*��&-�o)MhlO�S�F��M�y\ȆOH���hw \a�Ίg�ٙ���B��U�M�N+�`\}���'6�M;qi<�Kh���Э3�W��o&��|p�R㎭�{� �*�(�� ����2w�qH-��^�;��D̙�4$�q����HTx��ΜV�=�.`lM��26z�����/|A# ��� "h�d�G؈��}*��ٔ_=;^R�Dbr�8�O�}ʟ���]�(��!�Ġ^	ól��1	X� �͖fiP�ްZ��s9�:38�(��b��ݸ�zً��c�1EF�{k���f���B�T���������9O]���]�p�V�fD����:�Y�d:��u�.��;W��)��7IȉS	��K�ũØ��b�à�6�+'�X�&����ӛ���<�g���E%�6��"�.kB��D2И���Ry�����<��Bm8�F���F��X�a@G̍�Ͱg����{I��8�#�cV��%�`�Y�b*�g-�N�� �
�x���/�/�V��|�\򞊸S��GU���z�ړ��������+����S����vX�슋��B�ۅہ��T�)A�H�v]���J��=v�[�.�q(@5�ϟ޴�X�y|Ǽ�E��A�@��_�2'c
O����{<7��FOW���J��|���{��������Բ�b	SQ��js��s2b%T����ظ���~%2߾�k<��W�B�%���+,�5k��]G&ʈ|��Зq�p����6�C��H���LZ��LB���6����<U�b_��Q�]��3)>#ۿ����蒏��J��|X��5Sҩ�[��ރAojsꤌ��K�u�6L�k-O�?/)�T���Sd!Z�$*���?��-�d�f�!;k�(�p����U;}���������n�y��?{�(�Fr��SR
�\����q�t!18$6�|dO�Ϛ9ږ��Oj���W�t��;���qg�H��mxc�G2a��C�6��,����$7�վ_�8�1�=��� o8���7v�|s�ޓY���X�BN���B�ܳO]�6��+L���IĲ��*d�	��?/c��M��X�U��,�Dp�OhJ��-
�N����_%��N��4���X��|~�e�9���j�횲ױw�����`*������`�gݹ�����l9?E�����jʯ+$��.~8R����r99�~�jXV�=/!盆��Z�8e�h��Z@���|��FO#XS}o��B�\��G^���,�`�r�l��so5�
d�UlX.����Hc�ڧ�����V̈́?߀�+@��<�����NiJ�,Or�6)�h5Ǥ��L����!�թ0����������V}�擮�(U�]�dգqZ��h���c�9����1pE��|���r'(�+�J~���˺f���|�~Y9�z��Q����0b�[���l����R�P.(���~�1���<_�� ���$�Y7�a`�~(��ɸ����{Q�������(u�6����=��oQ���*�yq��f���F1���S#qm��f(f�*���흁���ҙZ#�\�X9H�P�����v�B���o�b���.�&��o�`�SX浤\�ϋ��WB�`"A�S��w;�1va�A��០��%��T24��]�ƚY8r�8W��&���cf�q\{�nߵU�c<��r��Y9s�yW��H��P��-iE'��@���C�M�>m־��V�#�ԱV8�����Lvv�jO=�2��crn�k����j��
|�=�t�].�	��*#d|��M��[ߢ�$�B�� +tp� 9���`�u;��ʵ�3ݙA�C��̍j�׍wt��(�
"�ḮG �>WJ�����7T�p�/pD�l׌3�Ǭj�Oq�ʹ��T}���[�h���HD&8�~6�C��Ed,�M1����x'�YC-�[t���\��;ZD��i@�W��x��9	u�p��`�Ģ��{^�W9�(X�န��(�o�+��c	�f2^�uKd�5G��U�u��j�$Fq7�BTg�")�C���C�24X1�����-��,�x��;Nx�1״�È�%�����k�
�,�ȹP�z.�O�W�g������
�����o���^נ=�YG�M�o��]��{�����F
��{���%�AqN�V����௷T� C@�65Q6KzǊG0$�m΂�a`=�8�pJ���5b���\��}X/+��a1���)��5�3�����!")��H
�*`�sG'�p��3�@ܑ����H��\�.�I��W������2�͵�^����y��~�C2�
0�NN�p)��q�k1����ˍ��p)�BQ7�R���Zu<�ì���ڋN׹{t6XJ�����0����� !�O$��ꔪݻ�8����Da���<[a&��6�ԍ�1�)������u�'z�2�<���2=�.�-�lrm��ٍP�I �F�s�Ļy8%)bS�w���Gة4k�S!'_g�]nbd%Е��Z�;1�s��j8���֙�ԧ�M�X5�Y��|�!���2"�ʺ���ixb<�I�N%�z�?��ƜJ.rr6�x�y�b�K�F#ɥ�S���&0�G�)o��b<sZĸ��i�ؚ�D���!J �~>�Y��aE},�Ƒ=՚��z����-v�{����\�����V���Y0čr�'P���|��7�עkg��.ج��%��"(a�x�]_&+}�xхǑZ={,� Ζ<�dhX�ㄛ��C��L�9��b. ��F��
'��rd����)'OLr�JK�ha�YjPZwYx���0�sN}9S�22t>Y�f�5)�(������LF�_(Ɣ�K���3\'S�p��c���A��Q����'H!`}_z3`���9�aô29B�w3DGaN�n�����vݚ4��f���6̧0�2��V�Xjr�;8�!�\�mlV�jL�g]�`�Ҷ��g�� �p����X�g�#*�{����_ʢaa3N�+a
K@��&dvo��o�j��b�����A{�އ�L���ء#ES0�;�8���`te�B�?�����+S�7�e"5/i^f�梘ǝ���A�f�#U�.Ƣ���ˆT�y7���/H�6���$Uu���X��|�W���ý('��:����G(��NèQ={�Fk��Y-��1G"�Ó�z�S�\�MO@��ћ��C�61�a?�W�a����(=2{�$1���e���:����]#����n��&��B���(�+D��2Q�vl�nᜨŋR뚣���2nJ�)� f1a�¸�fǦ�6t�OPYa� ���Q��[�.{�~s,�Q(�-��#��M��J\�X�h���)u������5c�}U���ܡ�8���!��k�	8:8�]@T4��)-�����4�N���@tiH��#�s���O����y�h\P�'����E�&�^��t�Mh��n7���B�le����FB�mMX�:�b�GR�rM0 ��*\l�N@�,��v�a5*\1Z�G�5t`4�yZ��M$3�DN���'lRW�R�o}߆�;Ž�9��rIX�������O��d0gf,ᇒ��3:_�#p���e2K�tڷY����1vr«p��r��%���Y�
��?o
���x$$�`�V�W��V�e�{6��Btd趐�K��Й|�B�̚>��F,rV$+�')�g�z�Xa��e�k�+=f��8rwvBGd��y�A��C/_	�{�����uY�k�g�h@|}*�l?�gc=P4-� ¼9r���h� ��0C����o8[[����4-P�Q�B#ڂYKu'��4��pq|�zIj��y�Y��&�y��iE!�4F�߬���������XƐ�G��0�k�DV�<�*��Kn�[p��A�d}n�G���򤮏�pUTd��Bn%�?m^`��@�V�|��oJ #,П�ݷ  ��,�X�.`��ǻ]�<�+w�B<�R��=sF�Zj:\+�=~�8N|0�#��mR�( �q�J�u�w��������[���_M����APt�/�*++1��i����K7l�N��}`(�m��&���� ��舘Z<�͚��y ��7��=f�\�$3$n�W�^���A�,��< ~�_&W0��m�]VP{�;��������Ϡw%��m�?4QN���ЭW�W1�[	��_�kj�1qK�z��OW̏��ğI/d�A1TN6�qY��;������x��%1��q��!�x���ux_cWR�Ƅ	*C"8���L��MTwƳm�Z,��nø���ln{P��v�l������*�E�e����K��v�{!~A���՜
r�h�˰֥13��W��b�s�&�����	���De6AT���2��i~'�I�mGM W�T���{G��� "�43����bo䐃��A޷���DεW�c�CYY�YV&�7=���@;�؉AA������(�5"{jKVɽ��Dś�4����n�3�x#�I��cW�/zM��Y�%��E$���Lύ^9�.x���[��+��b��Ɏ��sS4{|w@�A���~U� fW2@p��,����Xjd�Qt-S��E���[�?o
��^�T_ZL_v
�ʪ��$m7��E� Z�3�ʮ#�S��8�OC�r����l�U���vzT݆����|҈=m����$�B��a�g�[.9D�QҘ��\{>�A�©�ag��@5�R2�a�_����UN:1��9�e��oƼL��|{��vJ�p�*���Q�F�r������T-O��c�C���+^��.����Y�:�E���w�Q�f�Mf���������_{�1�f;��݉-L��L:O�d��k�pʛ$�s�r�t����G�]��9�g���-�;�BM�y�a/r��wy9�^�>j0�V�����b��I����d�xx�I��<���b0s����)W_[�C���p�C)����6-�6�$w0��s�1?qd1��;�ۤ�-{N�a�TƋ���5	��H\Y��r�x5{ݾb�!�\\*�=�i�I |�l�(�"]�UVsF(�Ede�����X)I�i�Ɓ�Ӽ�ߺ�߫�.ʠ�Җ�ܞ�1mB�E�3�O�X�bOS-�ցЧ�J�Wc>sݫ���Y�TϷġ����N��j.q"?�xbq���H��Q�{hq�.���
v8s�!'~��ʻ=u���?�sQ wg8�;N��ڊ_���`���@�޾=��W_�M�4�.�<��(�BV��tsM���~�Z'���4C�|.��O�=UԜ觜���cy@ F�3:][�ܢ�ђ��1>���JJ���z�-�
�	�,���q�
Qa���ד�Xzur���f��U��e��e�s"�g�s6+�e��~A;8,����4�䥧;}9��`K�d�Pb�䶋]��!�U"�U��oPS�%�A�z��X
ǳIـs������JbB�k?mb[W�� ѾS�c��XV?���)l;gh4�r�˙&��^7�s^=���G�ƀ��ާ�Ğrj���n�Z��<!�T8��ϨTv�K"��"ח�z���J+���ؗ��D<�ЦT�Y)BH�}�xL�9��?[�5�з%��N�{��:�;�*�Q�WlS���<>$�� g-�,I}�Y �
Y'��� 9��ѯ��L!ʖ·���k�����ïT
�� �8����u�L=�(�R�i6���)�헯�3Щ�=�g�ǧj��b��*Px�ZK!���xu.P>�YܸЧ�tn�f��a�+/�@��"KKY>gx�A<GQ��q�����Qu0ƥ�Rc�A������>͊Bp�l��t|���~�v ,,���-!�љ�hQ��'���
(Z����� �-�8ڡ+�!;+T���K)�E�겍�Vq ��t{����YX�/��.�@+5Q��e�,�'X�T��7�(���ՠ�8�n��%��j�������ԘB(�חz�w~�����ІRN5����h�()�GkrWe��~�0�>�8�Z�V?�c+�.�n1uٹ�Ǥ���g^�TO]G����O����o���������<�'^R2��ī:m�<��dz�y���M�:�<A�%#�\q�������Sz	�4�B��פ�͛��<T��N�SG�@���2�$�-����` � s|�jR��t�l6��֑$�n��d��i"	n9<��"�s�w�����iU��t&B���q��f�Пs���͒*+u����F�'���A�.(��9$^v��w"(�73��x�ʂ�eQN��3���$�T�aV�`�	�Z��{�m����������᎐v<�a�C�6X�{�����iپR�G�C�>��[���g7b�����hmn1H��"�;��9͙����Sl.��M*#��.Z���?�\,PN+�g�� �F�W�ni4�o�IU��w���{ʝLC:DvQ�N�pIz�����|d���T�x#�Lu
���y	��OKy����0�8�2^֙���_��#���[�ʛ��[�*8��"��0���1BWP��'��)�n�nb�]d>�|�"/�B���h��--�>�0TOtJ�7�yi�	�"(2-��H�����)��K�)TC��/��pf�f?*�PI���I)<Z	��ڹ8k1`E��;)9R#�9��n]��^xX�SSfH� DX�r�-�)��Q��[�c�!#���yE�\�ԫV�wb�X����!:�M��l����fʡ��'H��R:|��1��;�q�b>��PX���`/>7OA��X&�h7�޳ءFx�M�s~����N���EI�B��Z��x�G �������Z�(���A��$|��cU)�5��`J�Bk�x����`Gc�3t�4I���By,�cl}<���F��Ŕ?r��0��~�1�0$�%	*���Fv}H#u��=fjF4�Hip*��cS�9�vK4W�[Y�A�A��R���,���+�;hx�Cֺ0S�	 �q����ť�2k�E��<��7I,6F��x�?@�"Xb�9ΪUOˢ\�S�XhDAm��OQ�i�g��F��u���Χ�.yT��i��e �>^DK��Nv#*�S��?"E+�G��=��g�0uFp���,K��l)�ڧ�ú����Rg���2y^̲D-j��/���0$N I�{_[�n?�*c	 �er��g�ǟSH3�v��,�j(ͦ�C���@��7�ʵ�-=��	�*g�h[5&/�_�.eR�H�?��Q(^HX����N-�mhfM��ґ{Q����#U���5��پkr�����6�C?p�j����!�Tf���E�:�cf�5wv-�s�e1��sY,��o&��fw�>f�2u��0�d��l $��픱^������xaL]��?ց�it៹��<���%^@�K���9�<��	��O}�Wz;���%[G�V���0����2-���6-Sj~>�v���y�[���Y"Mjf�ͨ-�H��%�0b4�<q��Nڵ������ܻ=��y��ĳ=�ia��I��?|�Yv���|�؏�쎬��on��b�p7��Ƽ췠��ӳ�D��lK8��;�)�L/l^�3��]�C{YAw!��F�Ҧ�K7;�m%[��R�fGb�����C�j8+Kf���)�^��@�����=����7�z�����z� M�����z6I�T��ݜ�/�nd�C�$�ȃĎ����-.��3�4��I/ŠYw� �q-���T���3��<n`A��'d�l~�R��0uڠ���i��+f�0[�~�ߖ�#��O�pR۽�f��@k�`�z;i�<=����U��7�x�"̞�ECiֆ����;7ޔi�sP����*�����Y�=�8�I��3Z�b�B�p,=�B���j]�t���5�m�̭F��ƛUO��P��"ސn�|2{K���-����&�S�bB�Wv\�_~��.�|��
tcT�pO�� 2��
�� G��~�A#�5�����)���z���_?^>ri\�@������z*	���_�@��a�]L��l��G�)P99y�'].Z+�͎�I�z����ZD������A��C�J��0�m�;���YU����cv/���.��[�W���9nz-c�\���k���V��>fQ<:�6�y�aB�z"�%��js�ISU�F�ťG���Tuo�/� �LI3i�PHG#b˭�=2�
x
\�[]����yD�|�#BH�d4q���%KT�^u����8���F��f��@,l6�,�f�O����c��*��czt��o>F躌U�P��K����j�����Jp*Z�U�����9(�jC�QB����m��v����?�>Ş�[�:��׊��j��������$Ã7qKI|��?�ƌ�ĜdL��PM��nnR�is�t
�����XS�N7�{�����v"���q3���q(�Ī��v����n�~�U�tk���tV�]W��@�����5�	`�NY�Y<lw$Xt�ݭ'cnq�	�2c+wR���8c��E��,��T����l�e��C�j��D�Z��qb�V�[��&�'���|��W4�M�H	�?���S�U�L
�}C��}� �r�}�O�E���Lp�qx�Z	��m(w�G�ra�M�pD�M�4�z�$��y^��7�i='�t���bi�ZVDyiN���8&�4g�p�j/��x��~�{�������(�npUuƉ���p����fCi�A�cCۏX~=|,(��]��|BM-	Z���T��XaTd��n���N����	i�[ԓqcB��.�r��KJ(���e�Ɓ�&>����o�-�=��P�ei#	��KLQ�e�2���b9�>�Q��:6�N'��~�g�+�	h/�єI��Ѡ��I�^�;9
xT�JwF=�c��HI� G���*8{�iTJs��F��Mv�O���R��!���KcI�����_�Dd�$,����*�ʴ�\��a��K5p},ª���՗!~F�k[\n�<����Sf���f�t"�-)���4Q�Pi��f֒�7&[i����$nh��V0�mC��i���-+��<�!-`�d�2a��K=�r����;m��W�;x��_�`2'Fb�~����T�z}N?���"Kh�D�b7O��_���դ"y�����:~�z�;?d&zR��y�q�|�@� uq�+�Z�V E�����S�jd�m� ���	�5ݲ����nž��O�xf�|D%�����ϒ?��0���.Ѵ�w��&���(�Mi�.]��@C�Z:���F����}�2:�	E�&�j��I�jBA�^���&�,�*G�B��T���'w������T���M�ɟ�cbI2Z��?�^izt���k0�^I1?�Ioa��BMu[25Af�c�@@X�}%�pjҩH�-͟?a���\����WX�AE������dcsc_�[�XR��+�_'�l�;��8SW��H �&>/�����H������/��0p�����k�ƥ����m�S{��
;O�Z��~��3�+�dY���p #�ʍ�b?��<�ٕ(��M[��3�ƳAO\���Ee%��41�K�2_��5SoD�(aM��yW�=tRe��\Bݭ0\�U���|��$�=	�d�!���+�D���-,YP�;�m�� �� ������?+|��X�?���Z!SD����J�ν�ܸ3M�� �Y����6���=���z�̼�M	��Ns(f��V8Ot�l��Ϸv��g�̙��L2ӧ�_���|%��%��NH�{V��e_\��EȚ˥mZ9��;�Y�<-�koE���-jq��]�v�Rn��\��������-�jB�d=��(ėA�B�%,��̧(w� N��?K�F��r�KR���(�Q쎽aΉ-�O�U����Z�k�3�ʾ1�q�Vo�H,)ɶ�'Z�d�-�h������똒���W�d�� Τ�,HA#��raۧF�a�]�~�ސ�@��v@���*���ǀQ�X�Z�'}����k98�"%��R�SS�x�%�W+���b�����r6�d�J�	�!ۦC��au��~����r{>w���ά��󥻛_yU��/�8Qh���r�O�2�T0l.���;�y\H&��g��CP!r������621j� ������������~��'�� X���&�<��s��v��c>���=�=���pI�����/�8�\��r�~��ߺH�t����/���w�:РD�v����:߶AYH��h��f����
ﬢV�g��4j'�kZ��
�<�ƻ?]*����n˲4\��"q��� M.��j�t�=�mPO�"t�hP�X�� ��;"���.�6��wQx?���G]r��.��A���]	�U�+��g��E������w.꿇A^N������"o޶,��i 1�0���}�h�U�5�C��:��X��QDK3���OC	���?��O�*�{��1����<?�+ˡD)b�Z�c�{��<�rb� �)����M����P�x�C�z������i�<s���b^�=p.�^e&�y����b���;�:�9�T.��\���E��w���X�*i����ܑ���s��ZO;�OI��PŶ��N���T�H�uR�ZØvM���n�բ�g\�e�O�b	v,�M���`� ��-�B:+֥� /�����9Hvn�r�=�v_�c�`8�iDmL��\�i �ȷ�v9#>�o�[~�dfj@U��.�	Ѳi�b/�kg~�3WP�:��ӃL���^hb+�T��cЉ�H���e��䫈�p3�����;w�P�>L���f������;l*�o;f�_`�!��2�Jڋ��aU���_�E;��Z ���u�=�}���4��߸�+�Z��~�ɉ!9�R��7��
4�_���m�4�8���I��~ln�{x<E�{6B1�� �{W�䰝�!��/�ՙ�>��+���=���~�/��f���`XZQ�6��a�F�X��^,#F��\�qR�P����̞$\�d�,��"z�)L�	��g��e#�6��^��e?�I���}׮�,+Y�Ϳ�f��")y�.��5`���t`��B(U:� �����1�S�A��U��	�Y#mJ$�����F�P̉�Rp)���N�kI6H�;bܸS0%�a��՗�6�h=����,t����8��߄zuT�M'���^yʔ���:	���h�E������M�c��h�������~�Őn-Zb�;�"vY���|�܎�L�����'�k���Z�0^���#}��-�h�l�W�{�}���*m�*� �0��d��6���[����Y�{h����y&
̣�����S|��ٲn�:���vk�>{�!��)��`�Zo|J64�,�aE�Mx�w] ?Ǿ6eW���ktfl���4�ϖ����8{x������D�0�ۼ�t��oP�TI�E�t`�.w�it���/?�y�Kt� �˞�4�C�>�1��C�~u����
w�bB�$�S���fae$�:r�D=uS"Lz�C?R�I.��)d�����JF���t^��,y=~'�W+�=��åu��c�ܻ^�9�:sΓ$B�ǧӾ��ht��<%��9.�=L�	yUFMn;�=���@v�Bɷ�o
~S��~�ZO�d���$�%�w�{8$�b����g��m&)�(�p�e;@��|&QHn����@ۙ[��
�8�8a����Yb���J�#��G$%d�D�(���	���E^�`Ư7z���M���z�d1�{�������{|���r���=RH�������@9�.�!f n�,f��i�l��̫�je�6y:(}�ɔI-X�C��z�j�ju�W	��?��B�j�`}�]���,��������>��^�s�6]��&P��P��'�Dr�����9;H�&ä�`nܩ���6�\�˛��W���1S��A��q��z��n^�0����X!�3��,�����2-�����jE�*hC^S��dT���o0�R�@�"�q�����m�>n^�N���m�}�n#�CCȫAnH�T�����ى���C�����g>1�wd��e¡�G$}{��)����@�"
_��qm��z c ����uN�&ŰD��/�c��XI����pbn$J� ��3f�wGG��L�ݺ:/�jϴ^\���l؆����������Rf�u�bDM�������c�F� 2>��Hm���	L]r5���+�d��t�ю���h�Ժ���D�d��{H�D���L=~
�7�莀7�N�v#KMJn�~ $L��h�'����C���-h�U���
�7�@����ȡ���_��0�� �dTت�H�os)!�:�}S*��߬���h���X慫f�8~z��o�m�'��WCmu�hj¬ع́��	���"���4����f�q���nph�����]8Ə�����P��l�:<����/:O�\Q�e��U�%Ǭ�O�����B��-�:���V�J�Y�O��y�v�����Ͻ@�8Q�&Xd���V[Hd�4��<����,E��|��=���ӈ�� �Q�B:s�]�nqH'������}�5�A�mn45S"�uB7ǥ���F����E6��bv�]��ao�뽖��郣$(��>�Ο�ʑ2=q̳o���	�o��ߘ��#'LE����k1�6=q���mʹ�<SK�-����{k�};('s���:d�RA}��M�^�TX4�u1r���R7}s�YRj���5���`���`=FDDq��wE]�
�v|�ټ��AF�;�u�����T��c����\{���_�	eze�\��Z"έ[{\Ha�%t��vY��;�hXU>�� �`'��0ĮBC;6�e�iC����S>=*{3x"'��!��:�ߕ-ޟ�[�2?n��;m�x&M��/�����t�w��-�NL|�+Z��Y㇜�9����e������w����P�[0��·�d2蛖�Ot���j���T|Zf�R)��5��۟�}���̀{�8d���=�N<Y���Op�;�,������P�H��x��"��gVwS�P�"Q�c���p��k���!Zi:�+3�T�h��t��,Kq��]���1�\��3'�0��1����kc��u�>�n�����>���``PѢ��sq���D���$T�tw��R�P�OVd1x����=+u8hIĊ�(�����*	,/�k*}7�:���"���k�.-�a�95wyw��n}7����������r�֓+���6�!�E�u�rB��Zl�=�z܌���z�r�G������qk��!��'���e�g�]+�r���F_�m� �p�mz�ߪ<	��5�X�i��jD�I��SYT����T	+(�o�#�j�"�.c���I���
y��_�B�p��W�>��`tkk���.'9�`������}�3��b�D��0��G�2\�oў$�뿢�E4���t�7��]��
�?k���*NO�E�9=�P,"Ԅn��%�m���_�����7 j�����P��֐U���^g�V��4��=۔K6�fb�m<@�[�q���! �/1e�Q�<��z��V�7~S���x���7�>�i`�5�����!y�zCظl��*y�J.�Zu'�+�_�1�Q�\#:/���dZZ�1�l����đ�F �M�/&`�y��}|c��� ��>�@��W�N�/M1b�~��Z�ۿFQ.-g�7 |ђ O�Fq�D�>�����`^ct����ײ>	��s���@z��q�H(���qX^hD�O�}��M��Ƴ�&=���g���٤��<�[�bt��d�Tb�c~
�sZ�����;Osj�/S����"���Mz�=>��c��C�;&o�2;f7�z�q`�|LM���"+)�@�J�� �h��ϋ8G���_��2��Z�&��Ґ��
��@L+q�yy>��OӜ�n|F�c5H�PW|)��[Ƈ*L,�>��׍vZ��7����4k�bC�����t�/8�L��� �ܛ�g����;<�(��w��̼ZE~�r��q�1��h���/|��b��H"I��Q��p�/u��Ը��9�>��I�06jVB����E��o۰d܉��C���L�7��H.̫�I#�7v�kjS)I�\�+l��B��]*�}aA껗�V�]xmL�,����m8������`�`D1�p<>�{�W����4�
��h�O%͜�Xy_�l���$�R,L��'1��9*l��W��KV�bi���R�Ո�������ĵ'
"����H�<`g
�ߴ�2!�<p3�
ݴO�9�6����`8	��<��9�$�+�o_�x`���Lk���d![���GVY6���R�M� �?O&�b���sHHFk�x
l� �:�Q46��t���t&ɫ����bӳ-`�52���g!�����8����5�J&$?zl#!�`o�R�r��X��L��W���ߟ��l���2&"♉��א���;��CT.�]��o����o~�*�!D�^~?]�o@��.��JH�9�&��ԋ����:���y�Ģ�GP��l�D��3d�!u/%�=�7��H![�3%�Ĳ�tk8�z }W�L��9-w}��uk�u�e��J�`nb��Uԩ��U�B")D"uGL1���L��;	iJ���F뛏pL.xl2|�L5cD��Ì�]ئM��Er6%e˷�;�%�@3���5�d4FZy=�W��J��9�:��S��@'�/�k=^�jIH�/��y�ďR��U��Y��a�X��>N��&d>A�HDT��*�S����2|15�[�����>����J$��LR�&Ρ1et�lG2{���8Y���G�0zM�����P6�����.n��Z/R��x?�
Mܢ"5nf��02�u�p�ԅs�䳍���C@���ߙe�M��;C��4?�!��:��W: 7�TU,;a�����@I���c�c%;K��o��;�	�8�L#���b��E�A�ɾyp,D��J,��,����͓�|/��!C���f=��F���u�;��]���!�����\��Ǽ0W��K�QD�@����l����^��xP,:B�y�`�42��lQ&ɭ�?3�t�~�6�?�Ag��eR��Muf��p��K:��IW6!�v�\{6�;õ8��2�Q����`�Ɖ.�&�I�JX7� q]��3
����Z̟'q�EY]He�z��Y��g@���v�p��n./ق�F}�t;�J.�����^ �gC����|��B����_������-�8q��|��o-5���N���S���IKK�﬇A���-�	�t`ge'<�IV�(rz�	p5��]�^ج���ml��M�1� _�)\%�ӕog��B�aS�����'�#�w��
nc6�&p+-G�%G�������ui4fN&Q�8w�`B���I��d��������p뼵M����ka�����c���]�}����*y���>=�L��� ͒���n����ѿd����-�$cK��{�j)���^
��t(&���������^���|��}3o�� k������{��
��:=�M��&c�H��VD���5왶�Нi1	C��l�Le9�٣{��h���J݈��dD,�Q�7f ���y�x都����XᏳi�6
��e��a����ggy:/��<�������v��oK����)�����'�#��Y�_��2��Ļ���1ϕ��>�pP��$^2�]όs�<��s�h�\a� ������*��a�C��n�D�0!�t�i=�3�����7K���I�:��	�"`�(k��J���vQ�XW����Q�M��삎���@��4�W��ͷ| �u�	4��t���P���$e�yY��\x�9m`�e��q_���*nz�!
�{�`�;�����u�9�"y��=��k�S���)~�Ϯn����Ĭi�M�K�o�|�C3�F�.Q�|>#9F�^��C�ܜ(0���~I�wzҷ��X�6��E6�㡬���fR��k�ôy�6L�UVx�¸���w� `+e8`oD�̓X�7�cD�C�D�]�m$�ua�2�m��/�I&�Vz濴�2��b#�����A�;�7�N��l�3�.X�^�|Q��d���LS�{��b�L��9����՚fx���I;�n�}����m������ �'��ʂ�y�&i[�_���&�zX@~j���]>��~��o�2џz ��?�NmzKZ���Q�%|S���+l��'lx Px_}��]¼��	^� �����̳7��v��zޜ�^��l��Zngc��Ѫw/�K����l%	�*�ǒPa���1S�$m�h+�J6�5�z������sy�9��i�=�1��E��jf=sA�:f _�T�,~.)VQ��Qr�:_���� .�Y	4��J�)Ғ���h]R����i�jTy�σ�tB�����L��J����>x��*�/b�,o�N��E�� �qy�c�.S]�A��]���@�'�h�R�z��-2/X�-��� hr�[V��;��ԕ�`:\��+_���M�pE�M�"S4R�樔��!t���||׆^_5�����F�T�r�ً#!��l�S��J�o��Zv�|�o�s�V4���!���z��AN�M0D)Gn��ni�q�����M_Lt��d�E1��i ������W̏����c��e��ob4��iH�!��1H�6�IO9`y(`��jĴ��F�C����7��es�ֈ�1�l�L8jZ�?��9�q��k(uiG͓�L���VL�ߏ�a�/���r��^B�V���d�$
�\�X���8
h�ݭ/ʴ���0�? y��Y�v݇�jy��7!�s���h��0��ֲ7
C��E4:8�vy`�\��
)��}���D�����˅��Ұ�eX�oo'-�8j���� @Q�����e��?��@����� ����m�O������v	���z���&a�x.��"�����������:��W^���x���g��ɌX>]`� �Ұ%O�:�/���E�$*�H<��%��s	�����4bu���Fxj�t	��r���AԚ?����lB�ϓCub+��~X��e���|�yI}���c�7t-(I�g�7gx�w�oZ�+/M>��$��,�6wѓ�juKY���Jd�dS%�ں1�y�>�r3$f�X�4r�;f�z8�|M���.u8(�� hڃ��o��?�@�q���`�'�ű[�N��VX���]�ݗ�8}*�*o�\�3���2��U���x�F
͗�ZC�c��~4�+K��h=��l-�>�����"o�?j0 �p��m?�X'�p�U,"�I��p煘g�.v�\���@[�f����7��7	���)�kZm�ylobhPʠ[������/��>6����[����G��M���*��F�v�4���n4>�<C�c�{m�:�OA�˚=3������z�:ܗOJg���)C̏u��K���_Ub����K��(���' I�_��[]��)����+�Ex��/Ť�W��14z� ��L��3�jz�Cǻl�U9MS���Z����_Zu������Γ�2<�M���6Cpg�Ҷ�ڱp�܁�L�P~�BAf��o�!X�����zHxx�h�a�&�8lv��vC�)����(nb�t�`�B0m�dcl���Q�fbѩlk�gq
>����\�"{��˷U��o��c���u)O��u�e��6�R��	�e;���.����u��#U�K��-2J�ĒsK�(ML�D���������=���p��٫��_/38"������B0�橩0R ��8ɺ�,8u4�%�}j���nbL�|�c�Z�L˨�/��y)W��,C��߾�\�{��6���z;�2K'<��2Օޡ��/E�>���5#e��§P�=G�r��>f�x�qtO�X�ŇK8�nK�7e-�hQ��G+5���/;�	P)�.��^̣�
�O���=0�u�_ C�E�F��=��lSa>L��tš9Rn�l��o�2������x{���v7$\�-Կ�)n��T�=��@�l�"{h_�+<��pA�!�ǟ^:r�O�sa�/=������{h+�Ng�Yya�?u�i1c+�[�X�����	l7h�Eu#q嫐iﯻ���͜h����P�HA��ⶾ�X�Sz���I�(�yrB_��$;���`j�}j���V�Z�$�5օ��"��[�m}*�m��#�#U�3��*R¯M0)��9��j���nK�#p��˟^�։��
�I�i}Q�/�	3��k=�g�ʿS<N�J.::���q�|�c.��/�6�)J�	��$�л�gY{��Y��9L&h�Dm�RH��|2�5� �>ϬE��:�Hui�t������Ӹ��vG��m;N���{��D�8��.�E/jFF�p8qR~��2����&N;?���ѕE���GN�!"�nJ�{��!�I�̈́¨`����Q��x��Q�y���b�����6������䎝�^��!�1*0��bPSd�ʒι&?��H늲W��nڼ>N�:{�+�w+$|K�����x��[��8�6c�]���y�s��*�*ׅX�wA)R��aX)gn��ot���\�>�����%�_DBb�%Q���r�����w����	Ő�������
�jH�msT�� �x��x:x����,��F5b\C�@όG�nB=���;�[CH�	��Bvk�����LyzfW�P�2�Cj)�K���5��]D:Y1?-P�+��=�s�� �'�t��X=��4�e�s{w�����\ɞy����4��)lM�D�[��8�b��.y�TCt6���r�O:�����FO�3�ة�*�	k4�5ܤ�u؈1,���r�Z����xj�Z{�e�e�e�0�����@����~�G���*�.PX�%j�ȍ��
�6$k'.�I ț^�V�V9��IlA-��b��)M�x��~�� �wh}�nslf����Yّ�۔G�[Hø���/Gu��7#���{�����U�౉�/F�҇�=;��-.c��3me�����TZKsj3��C��H�������T�ǦŜ��j�](�й�wH�^�2��%>j�j�)-���e�bu`���ǐ�~
#��H�V�{��j'ou�cL�r3����
�(�^�w%a�|f�Hm.~�R���/~"f�K���-�L �����V��lb(p����TY���Rަ[t�'a��r�#�3��� ���t1T��8��y�:�̚�H�M���Hy	uߑcjkc+��]���}0M���%+�vQ@k~��AX�p_���ocq�6�hV7Q������FgZ�+h��KEG�$W�~Ķ��g��(�ƽ�e�*�E�������f�N�̇U{[�y/��3� �z��*�|4~�H]��kl�۝�_����ǌ��YM�&�ǲu� &��p����T����C���D)�<��ᡞ�ԕ�W�)8Y�(�� e}��]�O�p�����X�]��Ն�\������;)_�e~�<�J8�~����1����r�}����&(�h����l�	hz{����L�Osn��z�q^��}�Uo�V���f1*+nC��6�z��JG�a��#l*�h ���Y�Y�$YG�uBdp�$#~=9#/tI��� 	)��O[�~,Q�G��N�H!�"&6 �`�\ב�jT	�	�OVf��18��#䦗(bm�m�w^��?�sd��[}ϸ,�^�[]g�E�݃���I_�:NX�e�V�G�=�6�?&4	=o(���(%u�s�< l�+��졊�~���q�UؑZ�_4=a��R�a7�E��t�T<�%xe��tND���^=@�����K�z�&��u*O�0EN(C�Y����<2_
�ɮ�=a����Ƒ����4���� ߅�h�g�FK&b����u�I@&��� M޲P�g�YC��o����Z��K��a2�=-�!��^Bٺ}�c^�Z�H;����fp�Oܵ���gV��U���<I���D� +���ڮ��Y�5�Apؐo�U��6�
��B�.O(�ޒ�*�+��(j�,d֜́�Mf&�Q�+�SUNFjg2~-�8O�+~p��8�H��P��Ő���M�z��G�ޞ(9qU<���AA �1����ƀ�a�[��ך	�ݧ-G<G���r$����J"-X]�y�F���#ư�'I�D]	�d: ���a�1��J�#�ʳ�8���^봏a�O���MD�b�*e;g�Ѻn� ��H\`R��Q���"ݕ���~xf,i�K��Ir0�k?�6�O���W?�4�����P=P� ��}��cG��h;XBFb��8� ��%���QI���ތ�
hp�MEu�kVWB� 0R�-k����ѳ sB��<H���N^*(-�L�T;L$M�d-º�d
�ìy�v���G�R`���Ʌ48���Q��(��B�ER���y%3+���ޒ)T�H�/�7d���>%�[�fc88�T^��[]����3�ϼ������y^&>c��nO���q}�m�@�{��IÃ���]�5������r�=iV�ݱ�FH �\�����~j;q�p�X�0�!�׋�TQv�QF�L��u��w� ���u���ܛ�9d�`ؖ/e�ۙo��摣����X8�������s$Sk��t0qg��[�I���%�@,q�\� ���%4��	��ax�J^'\���P�E�?�ڝ��1��n�Qs�IE������ ��ÖJ�Y�.5Ѵ������e�\b��Y���A�d�7�
�$���,Q�/
�O�n^"��a`?i����0Ƃ0�.":�Or���W�6�n�ܡ+�0�U��T�+�e`N[� ����ViFwD����uv���|]��uP��K;�'�/u�����d�DP]�j��V'0�
J�W�T	�In��v_�
��&3��'Ɛ=�4R��ϒ����6l,]/�iE��X��.f� �|�~����ᬹ�kLVbΎ����,���wJˑ��Ӧ�b����������(��v��>��|�w�c��yx�f\*��y|�=sr��.��kI�C,��ot�̋�,ъ��\��Q��e)�a��冈�w��0�
�m�K@4�N;ӸTC|�ԅ�kW�׻�V˲;fr���+��9G�;��H���t|7�H�nz�*�Ӧҡ��5GTL�{+߭��y�q0���`"�{ނP}p�k�\�V��wu��M���3 H�d��H�K��kD�p�|�[:TA=��i�"^/N.�p�.:����is����i�����J]X�s�(^�f0 A#+Jlo�rG�!�I�ER��K�s�j��C��-�f���Qeu8��Zq�\~_li@V��Z�S�T�C�0z��Ώ�����	���55��v�l�j5�qi>��p��:
O����Д����DkUA%�y'�MZ�d�e��OQ�LyVr
%j�8�*G٥��J$�dR��Wx�4��l,g�U�-:��&zd�����a��Z�R#1(B�^�+F�3x�׹�e�E������U��y�d2��Ĳ:bGF�ވ�Ѡ�-���P���V��"����e[�m�=��۠OE97�)�\Y���w���!�WWs��HmpE���eCr�*M�$`F�쇜 g~o'E�Þ|~!��#O��������l��?�wFh��=��o�f�a�y��g�tNSD�ػD��A;c�D���GK�A�LQ�ب�<�ao��.���{���*�h�o\T�4��F�,R`yL���Z��`����cwKx�J�l@�=#�[���}
3ʌ�ko����E�\ �X;�ˤa�Dr[}�'ZU��:�,8�Cn�9�y�:�<���ʽN�q�hR+$넝(ۚb��Ԁ�fF���i����x��0�.�����Á�;��������N�JzOa%��ɍT^]��;[6f�b][�%u!*����8��1=�,k���jN�_0�'ڰ���廧��x���4���պ��Nq�$�wO������豟sá���T��fB����D1�t�Ql���r�$�×ZҞTSa�t�J��/�(:�Ȗf;��%Ͽ&���s��-|X@���T
f�*~��d<Ӑ&�s���54���9)�_�+�v��`��c��� �x/�n$Q=~,%���F8�St�z	ŏ�������'�a:�l&��[9��V|>`!�6R-}~$�4kd��c�y�UԽp-|��1���D�Vh,'x���e��+��Z�E�{�m�����.e��-N}�r�յd��LN.�k��*�hĔ/?H�����\���擦�ܱ"I���c���f��)�m��*��nxv��u۹ơ<*��3�p�C�X���'�xᓁЯ�Tjt�������o�,H.���H�X#ؑ���#'��j�lQPMm������;�{k0W�;�CE�&ylZw���d��	M�]H�I��{>d�k��x��U�L�O+��[����BE��-����a �	b��-Ȯ�[�^�w�XX?��[�� �]"��NQ�������|D�Ȍ7эJRh�V�؍�3��q�4�`')=�6m���2&�[2�+�E���$��}[>����0Hք}2޴�&_\d�)�w9U>=}l(�Cm)�Fy4?o�)��<N��G�yn,��2��|z��Xebw;�������o۪�[�o��	���Z�����RR��=��i��w�X
 ��l��)�vH�0�q������V�ħ_�S�]^�Aؔ�B�<+�e�S���(�U�|o��2g�z�9����
��]�>�?*W�/J���+\���$bx�����;
�;X����搗XHܩ5�d�!.��h�@�C�_,$I_��<��$4Kʘ����L�Rj�}�_� ��"�/us��3g7���G�� x�R��aq���%��U��SX� �n+c=�Z����k�|���n.����G��vF�0��z]�l@���"�0U\h�2wѶlHT$��H-\b�4�տ��B�;�/�A#脿S�p2��4�	%�wb�\ü_- 0P��}�E�҆���0�)�>���y��q1��?�A��N�<� �՚�7]�r�S@���Lo�5���Ü�8�Op7_ q��^E�l��^��9��d�7�>)�>����,]�ܨ�oq&n%�����~���?�`b�tmT �"�|�WLR"��T�F��l�O�0�j�"`�.OYk%���@������9��F�En��Cа�q}T�gQ�'\	���9�<�ƹ�� �������T�AvI\�@�K���!�m���崪]r��(8���V⋿��K�;՛:�3�ÜǮ��ա��ћt�	{�.c|-�,Eo��]1���]��F���G�Ԣ��������@,������d��75��	4��Olb�z�uL���k�~m��]��ٰ)�C�n���=��p�bz �n�=�wc��Ȃ�11�`1�<;��X�V���ÍC�?�u�oT�F�e��瘫����ssd��UH���3�I=1��(P�����fY�+��!�[*�u���KA�u=�ifBcj!lK,A�c��_��T��f�p<�l�J�n����F���V�#l�߇��d7�y�w5R��E�C�u�&�Co�h���B1�	�$��*���@��V�ku�+�������yo13��MbnRs����"��$�~F� �5��:҄��#�Uu�(�S? ��*UG�n��ꮣC��_u��H/�K������[�r�` o(=���v�����ߚj@�@�hw6%�t]�h�=@�ǚ�0��j��9��E�9t�h���ZP>/��Ԑ��M�W\O6n"_���Hn+���#5Pr���´�W�N�n�������ѫi 5$וɌ��/�Q�&����0��F8��0��ZU/\��xi)�!uFgj%��1%|B�H�8àK ��{�6�D4���0�z��K���R�Ct�߇�t�9�f��?�R-p�u;�|��z�$�m���-�#o*�gh_�+�i�1F���a,y(ٲt�B��TMb�]��YO��)#���\�0�:\��W��6�����,
������6U����mv���م�
��Z�B�ݍ�m�g�dH�zi5��R���<c�OF;�Z�:C���<68��� ��/
&%�~��ࢋ���3��-}��O�`�fkh��_2BeqE^NE���Xt8u���{�C=!�@�D�Τ�j��R�S�0���c=͏va6V,l���ɜ}��>F��y/S����?1���.��e�XL]�sD���s���?�L�b�q̇�L`���?��U���!?��`�D'~���(���|�n�;v4���+�FέG
��[lu:��Ӧ5R���RxIɲ+a�K>\��P��w�2Bq��9����m����5V����:��<F[����k>$H�,e��II��m�so�!U]w��J���Q4�f���-��⨫@@ �-��Q!��esQ�%���`$�������3(���?�(�,�/�(��`A>=�n�*b�sC0�`�V
H���7;LOB]��Ŷ�JG�ܪ��BAd�!f�?D��fR�>�в��*�s�dۺ��E������\\�C�R�:�m�,��G�-��R���5��hʌ�G���.����tZe�t�j/5~��?R�F���|nIM��ǅ����9�.��˛���Y������t;��?|
�4�&���j�֩�)�[����I�=l�����
!k܍l�⤿�a5��y�\g"�FA���T�\��Et�;�繶R��c�i����$�J���~{�_�a'�n��fdӲ�k���+��������\"-�f7H����7�!J[t�`&���|����D�pX�ϖi�����h��A�P&�QS�0��Y��B�n:�S�O�b�I -xpD�*��Gp�L����xr�r����g�����?���'�`�f�@7*Ÿޙ/"ree�(�j�W�o ��(G�Mʉ�{-���K��r.&�����O���G����̎�e�A�m�,�6�)�d"�����[AL~����8�0��ߓ�"rb9��O�=�w���(1�pyQ�TK؞>uL��[�)8�w>��17�jQ��N?�lъ5NΦ��~�'~�BcN�������C)�^���	�4�
���e���-��K��j[T^"��Y�t�'�N.D�{
Ԡ�� �<b`��V������P�m &��_���ż��f�-�{�/��Ai�s[�s�KW�1c�U��$��'���q��U�̅qazK�#�����c1_Xf-���݃rϨL!;-!%�;P
 � <�9T���2,W��O�-��_}�Y���:���o��n(�Ĥ���al�x!��"1t�шA/�cz����碷��*B�<L/m]�䳎�{��`%�5�1!��4y�4Ú��bx�FIKh�y�B�ą�7�/J��Y��wҒm����/S�9�V��\j��v�y�K�*�ޙ@s`	Tt+�E�b`}E_�Aږ���ka[ۋJxa\Zt>O��дp�#Ua�q����1�_�Tgj��{BLK���E�
�l��a�Ư��b�Y��87��M��ڎ9�����VE�xr������ّ��V߫tvo+z�5`fM����6jTg_��P1I@�����\�؞���$���_(�b�y���A\RJu��ێM�PD݂>��d�K����z�h��+8��Җ�ə��"�����%Sl�3���/Kg\1v4���޶�F#�^���~�C�:�x�x&��`,THm2OVҴڸ��͗wκDm�6�$i({��;kJ��l��ѱ�LVB�s���� ��hQ�c�t�������n5�w���J$p$��c@:�1v<)ﳓ%9T�.'��L=��z?[
z"�3X7����b2@�k�>s,�B�&	7-*Uc��,þ�}@��==;����C4\�߂"���st�D�n#�Ś~�'��x��7��~	Ы�����!��R��I�j���$��S�p'eo�(��v?���]�4�gɈ��P)�C뱽��'��4��Q���};��������
�\w�rv Tĵ�����Y��"$b��#��?9 ��_�c��=F�Fnx��F�Ҕ���V�g�=���,M�ŢN/cr��^����6�[�k"`*����+�}�&�v^A�=����ŭ�e���1��:dK(qjYR ����1mu@���k�DDZ�^��};�����NO(���t�D���>���>j��ۼ��M��_ks��G?�qE7���ض�ѣ0,u��E��Ļhv>`�<����Q��߷*���_�˨�L D�ʽ��gAĺM�$�`}�սu�����Ŀ×L��b�b��_R27���u����C�aXO��Mw:o����kW�~TN�W��B��e����,Ŀ�҅�A:t��aJ I{��ו���Iz�1���?j·O)��zhXцW��J�~��*��?�����f.��˫Т�{����ֳjD4Kv�E<sX8�" �K)�޾J(����7�� �,�X��o��~��O�J��2��۷'����_d@o��V%&�is(��z1�LN�e��]m� ��,wH'���Z�pލ�R�5�؊��m��B��j��C��M��3K��xp�Qӝ���V9��p�
f9h�C,�L�8�A�n��ǆ�d%}Q� �6)S����A�B�-=u!�F���.R2!��\d)u_E]�5BLY��	��_
�iW���6Ȋ����x�=��mtXւpXX�Դ�r&#F�KU��wDBR��Y��y�|m�o	6�2�!�6޵gw�����0��_�}O�I�HTI?pi�b�8>-8@���ߕ�JrFh�ˮʻ{����&��$#D����wv�7N�6��jr#�~p���8*�_�Ia�wE� ��*�[���!���5l��Z���O�;����	�$W�|U�\��{�'�STgL<�@�.O��k���jw�4-�����g�4�5kA��� �; ���v�и!��$��.��q|6hPA� i�z��)\��T�.��r90BF�S��3:G�saM�yܱKZP�bW8\h#�l=&=��P��*bwRĎ�wr3�%cP��.y��xd�E�e��f��u����r�����5���{�O���n(�}�}�� "K��f��`�_�'�k�d@f�?�Ap� e�d����\u�g�3�&]��`v��OLn��&��H��5z���66rEW$2#���/�}~����9J���6���#a�}�p#�����m$O�K��͋1�1����&iS=m,ܝSn�~�7�D|�o?���ߋAN�\m��k�j��Sr���>˴�{W�8���ߵ-�x{�/E�.,2�_w��\���co������a0�/��Z�0U�:8����a�>L�^��/��9e�BQ���Ƌ�2��x�%{�/�/2��y���*p%�����icu�V�9�_qQa1P����꾏���&B� �1k��d�ro�f�S�3�F��x��V��K���߈R�+0 "�yr�xK~>�+E�mRd�%�d]�ߗ��E��k��!���%��ށv7�xn)]�Izw�~�~ʉ��kۻq�!�^�� �H~^-���A���,ՠE ��Gn����ہ2��Qfہ6�ߵw��v�/��v�[�r���� ��#`,(ك��I$�(�~6�����==��+���U 1�uWjs-9aS퉍f�%z�M�r��s��{Wk�x�H�g��Z�oi�F����o*N��Đ�	t�!����Q��[_#$�V�6����&�����& �xu����W�Gݱ����<��֬oq>0DC&yg�Ek�_ۯ���:?� _�3��mb~*������m�������؀z`��p�A�3Q_[ۄ4��}�$��ݾ���V��z�R}�e�J�ߨo�I���[�^?�.������,C��WEK�%��/��0��>�1l������K�k�@��}0�&�7X�õD�;5Q�G#m�.�������p~D��-���������g5v�+j���Ck�i�tD[>����dl�ۜ&yd'�Zaިz!w�\���C%��ay �\�*k�v�p���cKu��5o
�q8����0Rڪ��h��+�Gf��=�\5\Y�ס���LIK�mz#"�<�<�������|A�(�<�t�H+���΅g��G��73��uq̙���'��:��䃇�}��������>�,ks�l�b��>�{nE��d���@���&��b�D4�ywEC\��(���֤��	:�V�虸�(א��/D�Q�,Vj2�&�K�,y��p�Ԛ,&=�|+�%Ǖ��P ����0i�j�tL���|�T��"=![���3�}�ʕ���e�p��	��z��2;y&w�Òa�,��7��Wߩ_V�NJ v�=�-�mVJS)�TUQa�嚳W��gw�Hm�C?�V��\*B�8*�m�$}$N�)�Zj���׿MZ�j�پ̈���Tۣ}_�0��͈�y���]�a+"��P����HIY(���;���,��	0@�"�)�p��9��۷�W˕�.N8U�����(8��!*�_OGAfy�;��*�9���"CqNʠZ8�p��:y�vx'��F�i>H��ى�a%�f�	 MH;����Il��+�u�k�3P��ѭ�����ia�J�%��M\��n��y>YLZN�-K�D��&&7�q$�6�L?��Qa� \�4y�����;�WU{C%�wN��g�v���� �fF���6��|�Laz?�g\��h��ɢ�ouɬ���;�qp�MP�[_����)S%�,�?3򼔶�u��MX�PXQ�N�:\NJ�K淌��\[��4��7���!(`�S������6I��/��[隟�r��e����o)Y��\є+A�)}���z�;ϻ�q1ߡ�@����1��@�ί�P�7��2ݐ�E8�8�G����J�>�Z"IMh�@��������x�ͼWb�:�~&r���#�G���v8[�d�'oX��i~
o������RGz4ތF��[����ñ�S�0M8���յ��{UNZ�c=9ن�K�ze\F��)C�y%ͬX(���PE2�[?y�n��}(w�/\�m:�5)G�!��L\�ט�x��I��s�{s��7�pT{2�XZ������,I����^�;�gg��7�l��n���C.���@�ip��_�h� 8�~�V�t�W���ː�l+P�"�����G��dK�gU�z�(�d~Ӽ����b.&�x��HX_t(u.���z��n����t+��m&K�؀W'TF
?1?�v����D.>��뤬��ò�H"�@0�ߣ�Iy�hV�������Ck˶�N���8D�ԑ����~��$��$�g�h�d�w�C�-R
�����Y�7S�[�ٵ�潖�z�*��#6�r�jں}&5�T���x�
U�$%@���c�̙#�Rk��hl2N�s����1$��_ �T���g/�J�	����,l�ؐkF���p��`���\ܹ�\���>�YWr�iuw�%��j"�H���F��&���[�8��+�	��A��a�ב���ٽ��i��ԣr%G�oU��kw�H��7��������m4h�M��n��׋��8�8�7�G����!�(���xa�i7��e ��8����yl��Ŗ}��f�'��Oslp���J�	-A��򗄐3g�}�wL��;�bi�¿'��Vs�������l���Ԁ" �Yz���@�������{;���s����6|�e?���,@l/��$���ǂy�F��$���8��w3�K8���'X*��`E����)VE�d�D��b��ۭ������v̅��2���.�R��A���܍T���1��^��$k|����8&����x� Q^+��LUh���+fD���#�Rw'�&[��i�#��\�o��b+��K
[1��teA�R׸*-Y��	.�2/ؙ.c6$Y��9�¡��!7���!��%]�-��X�}�o� I�^ײ�`�Htz�	�.�����I�%A�;��!4	�B �<f2A�U=��� ^�)�˵4f1m��Qr��B�M��NF=���RT��@*Im���M�R���ݪx��l��"%aB{#��{����\�	���/g��J�>	����$�-io���[v�5�B�4\MX0�$x-؆lH�L�i`N��3���܃���p�+�?�)�� &^;�j��\a��vw�$��]Hf~�F��r��ÊA:��G��
�|-W�z#��h4�S/��cK�aw'�̯9k�Ҕ��D�Z~%�P��y����ǭ���C��_}|��F�� h�hX�#ko�e~�Z��>Y��A�ݪA���Ua�.7P�.�t�8�n�8�J�ZO�
*N��SS����B�B�G��g�$��nΗ����>��@q�����ˋ^���)�M�#���ó��|����2cD
�pN�^^���Y���<�ǳQ���*'�t�peZ�����楿�`H o���(ЖE1���%b��#��Xhnrdpd�ʮP�ӯ9�?'��lQ;S����G��v�e���(`��Z�:*�M��߆���X�r���v��m%��֚�8J� �	i_�����h����j�z�Ȗ
[�S+?�_���!�)�)`���^5(�ˀ�
�j5��qr��wR"�������d�t��0a���4�X�*��A�x�A����\U.=��ӏț{����1)I��@�U'v6�3�A���ޒA'%:T��L����Bm���7<϶K3��H�.��FT7�E	�cb\V��M��i��L9�Ѩ3bu��.��H���<-Y�.��r��)��i0z����UeT��~�d��V����±�f�ҹ��+6�lw$�6�]� =	8ڒ[Q��n��#��M&�?�t�c�W� 	�����B��NK����ռ�۫�7~�)���1i��N��m$1��~����(ۧy�1�"�r�>G��XyӒ�Gq�������-�@��÷����³�ɰ���\j�)&�g�՜�����w���И-�D���N�]2h2H��N_���bz���CO83�* |����n���ޛ��s�2R^���i���4�!en!I��X�\P��yʃ��i�ׯ�r�9����U/)��Jn`?����-�#�V^A��f0�����$ԧk���H�;��6�VB{����B>�gV��ޘ^w|���u��x��)��� 0D����ɳ&pl?�׷f�G��/��)OOȻ\�d��H���bn���r�B�؇�@�����nQt�iK���F��,���mSu�;5agB"s��+z��Fh0\��B���'Ȇ��|��Q�'�K5�B��V�Q�{N�m���^j��3�UH%\��2(.w���'�
g�y�����Մ(��h-�'�ը=��+�6|$��`��h��ܰG�6f��>Qƫ9�d��&��m^ �j���XT��a%O���]r?�#�����k����~�Pn⾉���D���ec�o�6O�dY�t����3܃�O��n'~�AC�B�n��s����EGDc>��ya�e�����ύpu/�^��V ��c������W�uh���m�%��ˈ�����Ը�d���%�ǽ�9���$X�ڭK�U{IP���z��硅��}�f�*}����/PkO��f�̐����w �^
F�Z��4��HYY�U��y7j�م�"$ϰ��ˢ���1v�R~ �NR�]Ϛ?������ϕ���ҵ���e8Q��<P�]���2�oKB"�G-|۔���^ �<^O���T'��D�����b=<�&���*��"C�(L��ߩFߨ����M/CF@r�*l���6WHPN?�rtb�d-���T�T�eR)֯����&ʴ��:�s��
��;]������8b�R	�P�|���>SJ� �yV4h'�J��c���6���z`����A9#�T���$Mu��
\�5k�K
F*<s�?�Yk>�!'���6���6�jI��B~d[Ć䪇��W,7����/��+�A�E8�	�x�Qs$W67��_����p諷������|_3jC�<כ#-bX'*5�L�������Z�ml\�����,�p3 �2!SW�uL`�QzG�
��F��d�x} >L�b2~�hTl9xrSc-�D(��]�-�mc��,��&������,݄_re����j�_�Rl��>7]ȓ���X#ầ�z���G���7�:�M4&��ﴔ�[���K��A����`��V/��t�o��A��@��$�u�����)3w[)no�5Z�4p�H�z�@v�_G�)�X ο��:�b�%���|�WUwN
X����L�L�LB�O2r0�x���+���q�As|֊�K2��$�1�A9i��1�m|�C���^_��J:�s_�@k���i��$�a�i��ܵ��Kl�>�*(Z�r�^$|��Ḩ��
2k��Z	��{�h��Pq�S	t�,�������`�뉁��@������s��I�l0��:�>�o�R�Ft h�$��+��B�dg�gw�k������cp�����Bӎ"�� ڞ �G���5X�a�R���I��oA�]��"��qM��К���q�"����F��h�_Ъ�jđS#>���Ț|��l��KaM�ZH�k�
�)�!Ks�Hb�g?����rV�kc�|�<�%�����I��"��8��>�@j�b�áK�M�tm�y0	�T�C�q�'����:q�/&m~��:}��E�P�~$Y�:K�I��N�.ܫ����E����4��l=	ޘ���P}�H���~�S�
v�&LDK�|!���.�{$��5(K�s�����R��aJ�D ���^;̑V�W��bY.�s�Q9�1�'�|F[9s~��8�Ms�G�ۺ��Z QH��/*6� Ȣ�I�̏ǮT�`�1����ɵ9��o�[fM;~B�2ʀ�}�4|E��z+���9�j�M��N���������|��a�w,WH��Y*��b<[���8絔���-�}<�;N2!<j�-W�^
����6�A ��.X�o�g�ߒk�b���R��<��=[��T�$0�K�@�=�ʋ
����=�\V���<ɜ�`iK(��q�2��+��?
��%	��|���Q_6��K���E�%gϝ��ȗI���J���D��7�T0��}RX�����+N<V��u�PߪE�l��p^ȝ�R&�i�hp��[u�)�d�{�oǧt�~����ž�d7,GsF����Jwڮ/V�17��������k�$���1���Af�~�r��It�פ���iႦ^&�x{lwsP4�	�#$A�p<ۃǬ9�Y�Ǹ%�Q(p�?���#��s��r���e��tc։�,��e2F�_Y�o��Ѭ֓^�x7O�7th!�skR��#QX��#%'i�fC�v�g�VSXwq�>7�Q���<��4<;6��EP�GK��!I�֊�e~p��R���q��u�_|:�&u��Hs!����B������Fo���,����Ϳ��}��K/j��(f��u����U�5���A���Mg�n2��#x������ҋI^��zIN
E�##(p��I�w�^���s��j:���xK�>B��-��f�=ΰ��vh �b�v��G�Wkq�I!C�u� no�rc�~Mcn@��9�Un���V����S�E�a�{V��ՅaZ��M�λ�b�'T�}��յ�/W8A�@4*]~/�	qΏ̎��┓�Y[K�Q��>�����p����v7/����2���q�~���$��;�����ٞ�*��p%1{��b���zN�@�PV�8�S{UcI�C�6�,62b���P �w:ƫ����_�����F��X�=�CKs�L(�Z,{��uh�P@m�=ӆ %P��;�ݗ�Oo++l�-���j����ݓ�@��a`޴��FsO��j���ɲ,���v��S-���ng[�������B�dDK�~��ʶ>�?4�h���;ڏx���{�$��B_,'!���`ǼT�3�D��^�{���=N�o[�z6H㛂"�\�űL�m!31���>�e�55 ��C�ܭ�|�)�X�Q2Z��8�4Eq�<rޢo�6�McGz�)�����5Ӟ��"�Ot�8�������H%�j�t� Ak��.��I��׍}W�6o �i�)��� ]T��&�MjH��$[V�jlL/�C����$,�Mq�1;���Je��ZӒr�pS\�Y4�2�j3�V�P�8+�ߤ�U�x�
3�iU�(|��#��*�7��)Ñ���[�%�."	��p���TC"�q*��֪����*����V�tM������S�y`W<��)N����o�Ki��1�CG�@�$͋��@�l�3�V��NkK��C.�>�b��$�8�h�ѽv���lX��&�)��Ө�7��]��+���;G7�k��[�-^?���8��uw[u���xNt@��q;�� ����s��rap{�RQv]�~*���u���ܝ� ��Sa�ɛ��.�T!�F6h���Bޞ�y�~V��<�C�!x��9SY֒��J?C�NrW��â�n迧�o���M��uf���F�<,I:�A4�hG���>W",��t(yfh��,��tL��O�-w�T�J�,� �z��"��Ν~�u0�3_S���M��(wj[Y>��0afd���G����
/���A�1�������YV�Z�#�3��U���N����#d�c5|�ۻ"j��&E�����q�H�U�iI#��Y�5�H��b�7�.w�H�B&�������ڴ�T���>�准n
�(f��c�UyI�5�  DTF�d�n���ܹ4����2�bX�u��#��)���)�=���/�y�ʒ��ڇu�^��mP'm��0�'a\^G�9@3��;��X���e��B�Z�U�%�M��d�7��ь(Q}��u���xf�t�M�JO�5���^�	eѿ?U��+��*�}DOd��fɫ�`��Av�yi+
��a�TJ��e?l?���(S$�k���2�h���c�r��g�A%���g4[L��AV��8��2��7��dW�ާN�#��(�b���e+�eվ� �)p��Z�q;f&yg��h�v'�y�9��=q�k�X6���1 ZOW���h1��o�7."��В��"/3�`X���g͐�����x�+�,4��]3���ol^���A[��V>�`�o���4��x�]q�Q�7���_c=cA�q�=80�5䪬��h�{�=p�e�����Ѓ��%/t�ǂ��Gr8&Fh���"�Z6���E���j
�c���7Q������ֵ���q,�-� p�\��9 �I3���d�IO���Ӑ#%��s/}��ȑ�+͈%bXXt{����ڌͥ{˃�A4��B����	(�Z��+o5�O�PzX��
��}`D;�!G�;�G��H��S�6�m�)[��$|�Y�����6�xe���E�+�I�a-0́iq���'y��n��76D�^گrglT�2fGYi_ �4�襂����c�Ǐ����M�3�����
����ל^[z� a(���i���`ᕜ�S6�G1B�i�ה�@�4����Y�6'k���1�!=.��Et�|��"�Ժ�jL\�֐F�tn�����u;�j��k2Zc0��~����ʤ��t�c~�M�e�/�9	�*'ݽa���oy⭃���č`0HI9St(�RwV�US|n���`��j�n�NP�9`���o���/��ϋ�ͫ�ZB����E�@\���l��2o6i\�	��r1ٿ�_}ziVۢ�v]-=~21tZ6Z۬�y߻6խ��8x��8p���4��`K����)YE��wAO܊����q��V���y�2��}U�����NL���4���c��D�:1��QI��{�Y���i��օ��8�[��b�w���!��z0��ѩ�{�\��옕�f.�r�t�a>tz�o���4{��+��bx������h<��#P�_��Y֑dCvjO`f��̝���di��tg��:�j�J�ժd��Ț����C,lWz��JPJ���f#����!����.��~���j�f���E�����b��Ẹ���޹49t� d~-�1�
ܖ�m�?Ϛ�v�����m�9Jt��Mӝ�Q�si!{�h'���&ڋ�櫳�xϷ�n'[n��G�LT��p6�k,��(��=���d# LQ���O��t����Bt���9���?�/�����#���1F��dOs�@Ȗ�6��#F�AGa'�a�n������G1�i�̄)lvU��q�F3�.��)/�I7��2(��%��#Sx�76l�m��C�Ė"Wix���<�϶��h�͟���6G3��kvlB]W�s���bŴS�����wt	H����W�T��j��i�r ^��ATb�<��\�a������8�¿�,6����\O��>x��(�tꑬ���y&�8�����㓧�$*R9`йq�˴Қ)��]�q�sʁ��B6i����h"�����~*<|'��c#��_;N�ːB�����4�
�2[d%�E�^#�Gj�$7zQ{��	��@pF� ��y��Řӛ���Ҷ̗��x4�	�?S�&i|C��3,�\=�z*�*�7ǰ�Ǘ���1��n�|~��/ɒV��~�'C���{u���*���Җ9�9��1%B\��?���h��`�5Q�TJ^�6���d�	R��eݱ�)z�r�M�X�E��v�LQ����Gzqby�N�#��)�_fM��W�Ɂk�iI&9*|R��d�>S���
�lҁ���V���'��	\��'�3�ҋ��;�$�[)���/]v������"Χ��+��(��c����&�6���D�y��0Xaã�79<7&�piD?G�����+�:<��˝�����b��J����h~�ý>fo;���
l�ٮrC��^�����כ�Pj-�ε�<y^�L�9��W��ٮ��f��yK�Ms��gk����؎�3Zq:^!��*���k �a#��qFtcs��k��uy10��Ɏ�Q���?�VG�J2m2E�C$�-�����UWZA��6פ���6���_>]޺.&:���##%yk���"�=�<IM��Qv�!��i�����o�M�DC.��|e�G��#�|Ȼ� ]�����|IO7�%f]���U٩����D!��I��+H�])�sB����K����Q��h;�p�޳.��%�����`�;����e���������ز� �Ud�ԝr�!��JskeZ������4�@gΖ��I���9-,��g=�S3C��{� ͂�Fk3�@Kճ�v�Ɔ��^���iS�������9��s@��(=6����ݾ��n��ןW�V���D���3�<�F��ʡ��(EUHj�����E������
�����dV*L1��*���t	LT����P횜_�d�LA$��I#��1>����fm�O�҈(�d#B����󨥋7j����fG<1�W�TxD�����(Lp{�����G�,ѣ]�*M�e_@�1�2ƚP2�؅��z.�`ѽ�g��	K��8�.��Ӫ�����q�XRV[�w�^��ԥp���9Dy�Scx���p��eju�u�V߈f$�<�J����C�^\�o����4W
�m�值��F.@XEo�J:�����$��5h�����`(����.9��\55B�r"��F���7%��8��m���r)����%W��Bܺx��w%0Sm�����*s�8�G�^^�pV�h?�)j������Q�C�!�g�GA��p_b����_��x�2���{�T�����g���Ӏ��\�j�G��*�D�|X�{�'�!��Ė�2��˙����*��ω�Jm���4MӈpP0��[I(#u (�<�t_1�ƀ�aU?LX�gO�$m�%��h{FV#:�����1����ODP�.+�L?�f �,��V���}֍�7V��b�=�Ξ�|J�m�¬9�Oi��w��|� ��+��zX��R�O����ňܖ6¦+�7��� ��u�*6���`�y>���Mq9ʽ�7�ֽ��M����r-ˊV7d�)��y�I�e�T��j'���ő�`=�1�AO��8����B�j4/[D��{C�W:d��A���O�
t��"��i-6y����X�2E�.�5�� c;���I��źWq�������k��YG���̒��B�ϔT!?J�;q�{L�w��{{�[,$�y�^�"�w�D���i�ORFyN�Ey��k���]��* ��l�-�}�n}PM������u���h@�}M���+Ȏ��̪Px�ƹq�I�vc���&	G����Q=�*���QX{�SN�
�*����y�}��]����;(�qA����}�O΅ֲ������X
ů>�<.t��
��?���84X+E����k�l��%����Z@o�\e���1���&�@�����T�zz(c���Z��oԜ2�^gG�VHL��E��K��Ȫ�o��܏�����'ti�f��;�z���K�6�*?��{�ޙ
�_�����=a�fQ�|]U���8I`ԅ�Fu��|��mz�;ϵ�9g��p�G�S�I�VS���c�ˁteD1�v��U�r e�^䦫����=t7�o8Nv�Xۭ���Й1��uk���N6��To���I|� ݄t.�ɠ�]�O�#�{��~�\r��i�s[���b�0�W$�0�{�:�}d�+��а`c�3b3��s��F!��M��R�0�PZ����]'�p���\7��L�q�#���_)>��4Up^�l�Tf�(���_ۂ��-�z�"{���~�c1uZ��G����]�z6�][N�J>�ə���)�#��c��D���z��P|ͺԬ�����6�x	����)rQ��R����:�CG�y�c͔e�c��u��0)��B�M��W�}�{$uv<����%�/�%bO23Yci�Gگ飦��6=Y���7��<:@�Mlj>@O:́���:�X=�pQ+"�� B�1qh����c�����|)�GZ���Z�ћׂJ�a���/T�턨�g�>��q=)���j�a�������Z���`q��������2��D�E=��eA
���Ju��o�;HT.�$h9>�n���/a��NG�#�"�D�U��g���i,���C��B(W�Qyx�CZp�м�|q���SÂ��D�rN"P�p��Ku.6�Ÿ��s�:�e��h��F4zGƼ�UcK�U���n2��ű@��']B�^�(���S��Y���R �za�%���w�2��܎<a�jW:J��M�Z%�?x4U0�pm# �Ξ���kU��O��K�T�o4�xY��Z��j�@N�1w��O���bq��(HL��ϟVxкY�M��c�����<=?;T.�����2p>��&�7���7�"�����@�<� ظ+A��,Yf���+[\	����̄B2��2j$�;����>d���<>�E�Ɯv��C�v=e>N��C �������l�W',�@^"t��ށl�F&,P�������yx��~��:i�ס?\��<7��X�A�8`��g�x~^O �5,䉿�X�V� .>}8IA_i�e�h����@R���V�8���B(�jϿ��v(e@X%�(L�J[�סA�f�sn���m��k�"Q��G���P� ��oQԂgn7��@�bn��1=�E.B�:/3E�w��8A��2������2��3)��m�84�����u{��-�U�������^��n�#�"ݿ�@��@��<�7�I��.;&�g��@˯ "�1.,�}h�"b�o����A��>]��n�Fv�(����Ò�̶S�8���\���� !{��1[�9^�f�BT��7�c������H� h���^u�o�%���ś�0�1���N�d��.��k�`��l�b��3�7��1��>4 ʷKwft�l:�g����Oev�w�@��_eD���q"��n�9��Ĕ�m��v�گIdGb�L]o/�kr�k��u�
	����zT������<:��!�17˞�p�+Zv��%��
1��-^5�o��1?�'��(M"֚�)WE�M; Dcľ��#B�E'�UϏi�ʉA�֏�%{�T�P�밤��O�ac�\jҩ)�2 �ETX����m������Bi*ζ�ׅ��Ӎ���N �Z�%'�)V�a��
ks��0�������K(U��ۼ؜�Cu�M�'�*`S��aV����57�H�g-��1�����x�DXxW�h �nZ�s�B�[hGI��%���9�i�,/"��f[�P��`����:M�Ћ��aiߥ�c_u֠Z"N��4Ⱦ!כ��=ą��pה�Д,����[�3iT7�=����g2�ui^W�t?��\y��t���,���� �E쎨��tXݒ>a�J-~����E!+����1�k��.ჳ�RE�a�7��J�+�2��o�#�pT��7��k(�����j;���pE��v-����e,��t�C��d��<@qv�qX�z/�&8�B y����̇J�B~$ς �l_a@d&xzt��B�A�$��g��6�a���A��~�*,�j���/#a�j�G�|  ���)7�,G���BY�LNZ����%���O��^�N
6���z�s���aYs�d�`V��`)��F�^8�Y�9b�k�5D�oa|��v�ci!�
n�fB��EU�OS-	��+bR����+��5�J
2�4�ѡ��U��a�t�I�G��)�f�Hwr�_r8ٞh|�#9�bwCF���N���Ux�>����ü��H�����|5����#Ya{8{.��<"�.��2�	t��p^�[�SZR�#�q,�w�}<�5=�/+�����-1X��#��=C��q�����Ӆz��C�㽦o������Ńk�#7p�
vD� @V �	�C������_'�OWgj���BN�e��kwv;t̘MC���C��"��a��H�29�W,�{��?�D����0�r@�q�i8C�b�]�<���&T)���E�e7��ƍ�����g��h�@w������)��@�Ξ���\�7�c�^`x�h�W��0g��H{��S�M��?[��>���E�Ų��$�moƣ�%�ٿ	dR]3�;p���)�l̐�k�94���ԥr���l�n��{
��HT������M\o��O)1��#�Mm��W��_�$���Ɠ����B[��46��|����/��y���g/��N�`�h�^ё�g��k}Z�t�Ą�MtE�K���h7�d��^���i	���hˮn�)�=V紛�5��5�`�������W3e3>�rH;ZQ��ۖ�q��Ї[E�dOw�p]����{i��c	u�0F64kC�)W&L�x9�|�����2�j���Sٳ��>ԛ8t���q�Uң"��<wsK3`H�˳[D�K޾��vk����)tC��L��K-��xc�c-�$��lR�ϔ`]�W���ӟmU�Rޜ�����n>2</]) B}g������O>�`�d�$ސ���b���M�MQ�bBzd���$�"ﭟL��WӋ�{��G��p{�L8��o7V�[���M��'��=QV�$3���F|Z8���K�}(G�P�2���=Ͽ�|�;'�x��F�o]�^J����H⿚d������^
~#-��SaO�È���	~��Q����J�����1!�b��]�hf#���<;����I����
IP&�J����n�}낽�P�Ě�%�ZC=�,&�����$�g?����O�F�)a��T�t�� �_B+�k���  q#.�k%���)?��d}�6���O�uO�fZ��5H,�h�E���&��CҞ����M�|Lzi�ɗN'B��Ѝ���*�������L{�w�_;<,䗚�R�vP�5��XֺY�n`�yfN+��V���~eт����j�����\]�8hb�ۖ�;�K<M29�͙Ǡ�8����4q���K�NV���?i	tGO~��n���IkS6IƆ�(N�x�~^SDr�nxcf7�n��f���Ϭ�4\�VR4�Nƿe9+�	��&�oW⁦G(n��f)� �6�
���e ssE�z*�1�����>�dH���B E6?RG}Ƹ's�-󖿄��1��U�_��b��
��x�j��j�����9���~Y�`����j	+,$1}J)�3�q;��ܓ{����UQ�[�U}�V!������J�T#w:����hW��h2N@U.�L��7ͩ�����A�Dr��[8%cE�ƪ��A����/=�cQ����-�S3�5/?��q��b�\X�;��O\�q�x%�3e<��y��Q�UR�xvM'f1�2 6���{�)�q2:���� �Ę�_.TQ�X��_�΍�􉣳0 _F�]��\`<vce�A�Va�P������d��B�bP��3a+��Z����/]��?��wq���>7���`YV�:�����ĭ�A(L����,Mj���>o���GꌒcO���J	�������9�5��|V`���w���|�!�)����`�&�k5�Y�g��4-��r��@�'7����Y���8����@A�^��8��/ 8����o�h��=~[�t�����sȈ`1LC�g��xn��`J�o����W��C5K\3�e4,/��q�gg%��R#Ah����4B2���Ǘ�y~A(Wɡw�u�����tb�n��
-�J����*0�B�kMn���9_r�ep�+�<�Bc���C_��j�0ȕ�d���D�<%>��^e�J�~#BD ��\���i���7vw�����|H��P�bW�}����{m�J����LL���ܳ�5j�<|gή}���8��\��(?P�D�������F���[�����V�;�`��z�0��.n]q�	dT¾ v�;��j4?d��ͣ5�.�T�?6�J���T��ϫw�'��a<��EW��ft�و��)�Y]A�)K�����+}��P�W�/��Lw����8��^�H�}[a��h ,f{�V�̉iNm��<?{u�du-W��r�臬�	\��Ha��u���}ӷһ�	J�k֧���^�:��6A��MB\� �����x�`�/�7u�[��$_E�b#��;����	k��.��}�j�CB�	).��GR��P�f�c��,->=�ĩ�'�T�Ⱦ�H�B���!4w����}�_q��^��CU|�O�X�Ts�$5ᚯ�7[��*�KG*�`~���/4�a]��?!�q������j�p$�����,z	��
���F��9�MC�,�t�#4����4W������o�h�7�-�4*��WPds���6�׃�cB> ��W�8
]�6��/���:�"�s�E�1�صṪ%mթ:-�3Ȉ3VKǒ��P�	��� ��bg�0�y���gK�;�m�̇Xa��4�NR���u���Mb%��$oҬ%��Ǐ�NZ���`S#CT�[����ޡz�WZ�7	+�����ovJY�~�&���?��������撬>�i&�F�wG�Ě"�G%��c67?�/�1�=l�/�����5�)���w{���}��Y8;���y<aÅHHZZ� �2�^����ض��y.�����H��KV+��V�T���g��ҰG;�����N�.p�E�qe���!�!�x߲�ް\�7?���H\J!�s�Ʈ�
���6�fdEz�s��qz��G�pw^����$����e*���T�#U�c�O�@���x7��W~�њ��C�s�iuU�zy��p|������Z��sG���= t��g	W!�*��Z.�hA6�������C��kp"8�t�)��ʬVxAN;��6�3�'�J:�5w�`ٜ���t����ޥ��=׌����GAX ������O7d�=7`;�.q�V��G���ru����މ'$����k<l�ɢ���9t�{��6vv�Ŀ�t
G0z4��X!9�z�?�Җ�C��u�!����PDϑ�5IRDq����]����!���&��b�<J:�����S�y��i�~�5F)���CK�ѿ��8Z�f��C��l$���g0�7�m���r5�-��X�q�C2�\�3/�:,������@��HSO-n��B�"�����״�|�%��aPY��n bXr�}@�;��,(l����ma{���ê�B�cr�����"�2��6�%<�@]�D]j;�4��I�&o�崃��x��=^�����79x�>��fR��9�Y��$�²�G�u����1u�O� 알56�;�GV1=�42"�[�o�j���&j�:�e��B+�4k	�v~
|E-�o���[�����Y1EF`m��4� �dF�L6�hr��Û��b=r��9΂�&Z�7?�d(�rB�m#6��஖���\�:��Z!9e45<V3�G�5�@�L`���9����`���pK(���5֨���U_]�S{���ž6D�Vh+.���;���)ۘ\�;5/D�����ݵo4�3m��t[���J���-.U9��'ښ���&?�w��)+(���u�h�} �	2�eU̕'@�@`�ldJ~�~i��#?��ݧ�p���]���`W1�v�=2��貞������UJ?� �[?_]Up��"���#�	�k[1*�H	4[s�?�J�-e�x�aQ�x+C�6���{�9�����U~��s(�P�O��Xp��ϒ�/��ZPET�<�T(`�@���v8����i���V����C�F;QK�#���o"M�r@-��B��%T�=%
��ygέ�d�9!�Gڠ�8�LS��qwa����>%�j��6d�(
��VȻ����zˆvʋ����&���>�]��.����!�X�Tvy֜y��9k���li�]㘿�^��b�����ߘA7h�OM�X��֡�V~�y�����7�D9a+B)�
�ܴ��7�y6Ru���JX����y+߁Eh�ߌj1|I0Bh J����?Un�q��	������;+�����M��낺h�:����(�������.{���J�.^ό��Biو t�����-R"��YbF�^�9祖���R$�]�XM�3<=��m�HW=��P�mxO�#v;E^\�����<��{�*Ų��^	6��ǲ��G�����m�Xf ��l@D1d���d��H~�gX�B
>(�}���[�T�	3���D�=Q=����J�Q�2y����_5�� ��`3�P���}�&(r��r;m�ۅ�k�j����P\j���(����y7�r@W1 i�V3�k��OU�|�z=n����;w]+�0��s�����#��<D���O�%���ֵ���o�HP�ߙ���PB�a����� ZXU�,a#���a8 �i�OE�b
��d%#���0b�z!X�~�D����U��F�`�CY�kx\o_����o��D
}a�0��?��2�Q�{�)��>����%���FSa�,3���6p�o�-���2+O�ħg]�̒gll��Y��܌�0\���~y�P��PtAj Yd�cUl�0�lPUR�0S�B!�"�����ٵc�է�G!�/�b��FA���W�:��PX%Xs��#w���J��:b�pf=mˡ�����C�T������2q	�?v�cO��` ���g>�*tE�:G�BUv���:�q#	�ep`]��#��yg�L�_����6	�;���Had#���U?q1ᬏH��C	��Mu�_!s���x�5��L&
)�������&W!�#��� ƫr���9��~gWg��A~�(u�<��sQnH�̝�|k�T�LЬz��J�]y�j���'&{�>߭�GC�nM�C'@�c���z��9��ݥ3�g��B��� M�j�ki�\���ʋp��f�^N��z裊�ܡ����@n�UR5򠬈�A�}0��ka�����kԁ���Ɓ���f��]���ݍ��í�6 �Q�NyY�0�K�p�k,\C��%@0���\z��6b�d�e4R4��U��'S���޾:���q���9�>��#�5�9X���m�¬V��+����'9�s��8`S,�/��&�rQ�{��q���I�5���?�|]z/L�[�7�w
���\�Ux��yKI�э��z�_ H%l��EA�	�k��x:�85��V���M$�f
��[�Kv�d������'�C���ݴ
� ���on��f�����$g�
v�jz�	�F�w�f*ӭ����O������=H|)C��Nm�ڊ�)��L-i��2�Y�jci���!��J|�v*��k���s��o
��F��V�h�t6]~6��,��5. �=��x�)��8�����I�� y�m�7
qa植����K��E ͉ս�Z�YW�Bi��/'�~��>��T��=l�>�_`QM�`�3X$��6��y?8���<��gy1�T.Xhm�S�lxZ:A���p�X��T$%��m����w�������ŴL����C�Rn<�eIM�7��^?�1E���Woܶ��i#Pړrm{"Wr���l��u�ݏW�w�N@I�&fa����q�9�4]�5� w�xt)�uc%/	n��[�pt�gt�|�z;�)Z���t�kD���������` ����B�:�}��<�%��<�T��͇uG���'�pg��A7��v1GV���"
H�~)�+�"�����~+c-�jQ�]�"j���x�ȗ���=�t0�F�`�d�YFƍJ�]�UL� ��;�H�T;��yF�5@f���Z��ð(��Y���לXs���*��9���x�Z��_������ٱ"ʁ�n�T�0!l$��VW�Z�c���,������TL1]a����l��G�	��d��a��W��E���%t��I��<�6E𙼫ؠ��|�y���S�>nE,��\j-ؠ������vω5Q���(�۾���'�1o'\z{���;�?p� ,{-��by��T�6�<vl��XX�/��gC��=�2˫�{ң��!.F"&	�Hp�ӕ�|��'��!��"+e�p�R��|_���JWc��!��a0PgV)l%IU��O��=�N�\�k�2�3Q^����Q1?���p��I��h
�>OV������A��_Za]
�m4�7�ô�ī�a�OeJ~6A�I�_��7�C2�BL|����i��"J�����bK�V��]�/n���� �������J���*q�.��U�E�gZ�`��J����!�?3��Z��M{"��f�����IMؤ6�p���O��dU§�آ��N���=�r�hp�M�θ�͸�c���p�VcS�|�G֣��a����Z$g&u�>)�t�\�U1`�(��.Zi�R	9��dU��񁛈>TGW�ٍ�&2*�Ϧ���n��S�(��P������F��"���07q���\�v�J!ĝ\ˀ\�oݷLh�E(���5�{�><�%��(�9	%?����?�dW_x��K5u*Ӝ�f�*"�ݕr�c�z�H]��E*&5�,G�``�q	����97I����[�a�1��:����UtS��R���P��V�
�G2��&x�uJ�w��_`��tl��7�=3���9-�;���v4�'�����&�zK`�����C�����3Iv+��	���g��&%��rgQA�0�q� ky��*%�ݧ= �JY&*��zlD����	Z���1��<G��V��<�s�A;<)Ot�)�(]l���N/E����ΘL�H�F;x~���ϣz�j�{"ȭH���Â��bp����pAg�z1&c����6�GV�4ә�>���8�\���°�CV������v��.�N��d ک�m%�~Z�ݭGI3��RF\�&�S)ZUZ�%��V�M���������oaN-G�l�DG�h��,ڬ��Qkou4���;�[	��K/)�k:���2�ӯ*��}I�r#ݎA^3;�:*�R��#�?7Lé�[ۄ�QD�����Q�
p̷t�L5n�����B&�P@�Al�0��ej���nʿ �&d����� f��
iM�tY��UJ板���9��Kٴs8О�SO2�ҐǤXB�R��K��[L|�\JE���<�I2��{�3�K��P�n����T�����w�8L�G
��į�h��x�H��)�j��C��T?��s,׀��B��Ү��`�Հc�f��W3;���i(l�p�h-��6c�PU��w�ӨH�36�׍�Y�[�����1F���fʉ9r�E�P�be㩢�dUj�c3ZNmF�����i�Ug�3/��o���T~���Ƿ���_8�Ä��md
S���x�������v�+_�g;�� ���K��a}�)l�����e��/)��%o��E���veb`mF�t!	R�ī�"K�����2���ј����PTq�j97w��B,�,󙊬`�O+���JP���Ģ5�x!��'���r���,ұ�1pI�Ĥn,��YMU�¹��?���R[lP�P�z:;���p�v��U�%
-�4��3������l���q����pܼRp�NƕHLIR�p�=#��ѡl�`wxX.�^����������_��;��7GV
��L�0myI9\pc$�˻�q�)}���D ��)})�i삲Dj�|;�u-��d���0�Ȇ-.ޫ��Z�d���1��+�YXx+��3�-�+���sEm"��I}i�#�|�� ���t�+���$7���6b[�� b�#yZ���~��#L!�3a�=U�}2�<j�N"!�j7�j����(k>� ۪�p�&�	kӛ�'����,{O��6��37�xhK-!K�8?v꘸��ąc���#���(�d�h6�<���5�ʧ+��X=.d�W����qe�-��m����h��CϿHu�yi�oT���˕����M6���	0�4U�eΞ�Y[��-r$�l�I�Z\�̴;�=CQ��)��"t�<&d��T����_zg\��3�'��ꟳ-�ʼ$1)-;y�d깓�V�k%��V�LE��d�'}��1Q���|�^�G�d¿zf���!��}�h=k�������#Q�K��4�ϒ&��J}�_��X�D��3l�CƏ��F��M�����c�u�:J`e�?�Jy�j��R@A��$L��/����z����-^4�3U�j="�+V��NV��ݙt��q�������� ���'�Uz�����s�R(�rY�'<�lh��s�[���s�H��]�X�vH�� ��Cx)�	_��G�P)$f����.��69�n5]��G��<�?�L��Y��k��+.}�1r!���U��	 ����j靼t�}�r�7&����&Z5�9���:o����B)z_Hu��t�s�1�6��E�6V:�c��.�?#N*��,]40���#�
%6`j�p����Bw�pɸ�A��y	�'K��=*��扂Vƫ�`0`'��w�Ru��L!����Tg�.a��)��ē2x���:�ڶ?]�J�>�>P���i����A�٢�xO-���.��Y��_�r�BFq����L��YTMR ���_���*�o��®]��\���>�b_��+F�A��+�8�2�t�>��<��?����
��ڡ�����-V��L��-3a�C��� �ؠg�®?������'�]�����7���_������|������*�����7�P��p��K	<���eΈ���Mw�H������ErgF	���!��=��BF:A�9$���?i-{&;,�w�|">e�ӽ�a����b��s%I������+��F5�U	?	�;��x\)�0j��|���ӜCu������b,�=R"��mX�,[���Mz�k�!���Ȳ�{nqy�	m�StԐ�%��R���sYt���)BZ�]K�j5@D{�G��,CKG,��9�Ehq �˔���?,�~��>����.PQ�*?X���9b�k���a�Z�eD[���x��{�=P�F/��Նa~�@�HͶSE�e�߻� U�{�e��B�bP�_Ȥ��Z�z��B��oÏ���`�&��E暭��krֲ^���#�bqJ�F�4��W�r��^ݗKƋ(�������v�_Xof��f�����j}k���Z��Lv�x�n�<��QDv�^��n�@[S��[9x�g��k��/�5'D�'�3�0'nhU���6�5��,u��d62כ �6��$�8���I}ә���~��T"�N8�Z%���Ǌ|��\�}?��8ފƙ�͍�yX+�(���$���Z�D�n�;�/Y(�y����G�N�k)�rL�J%ߛI�q��z1��\(�T=6
�?�����2�����U "�����e�4�iQ	S
�S��FW�u�u%�������K�о�T(�D���A�������VU���$y	2\%Y��%�$с���)TR���/�����d$|��Ū�^��#��[��aɿB��e�v,��|�n!��<b.�S��j�V��Q�M.S����p� ��K[bo����"�].�tXx#�7R�Mˉ�q��K;�����x<麃���������KDVg��uTm[��2��ǜ� ZyR0������z8V����֜�����h3!Q���]@<�,�Ә�&ަ�I�S/��(V��Qπ�Q�6{�R!�೑+M%���A�Z�e��t-��#�����L�Vli�Y�i��L�`�TO���@�?��S߫�h��LN���D��F��t������'*�|���L ����θί�M,�[�t�'��=v~Oa%qs4�PC��R�3��@rq���ä�?��ƛl�\��[ G.=��2Ǯ����v���-eɧ-����O�Ϭ`h �9�0N�7��0�����y%:�2�..j������TO�U��y[���AGa�q.�c��g�
:\	��n���e.�������T�a��T���xO�����aVw�2���N�^n������+�Rc�ýE��\=x���Fl�J�Z	L^?����ɴg|9c�a��w�_
��6�u)�f�t*���,?�=b��[�Xs+r>]R���-#�M��#�L�����	&�~��Ģ��v�[3�
W߽� ����)4�ꃇ��oF~���ɭ�����=��{hP��4�8S���
�`ӓ)��V}�$�6*���i��C�+A��F�w��c����b�j�eܐ!L��:$�
�]�v^��Mg�Z�|�+�����Ր��H�$��f'��L�>ig�󑾟+4/�?ޢ��l���2d#|�Ĵ���`ʸJ]�%Y�5�6;쇗%��R�N\�\�D��숺��Ӑ�`J�A��x�&��r�:	m��,=���q�lٻ�L
2t��ܚ]ܕTi��piu��@��
+� T�b[`~�ᥩ�ehܱ05�"[5���2�TwQ�d{U(��L��\���l���n&ꡔ���9S�J�~P�� L�FZ.�~!T�����/��e?�|�I�'�����1�!n�s�/�V��d�?[���YE�ǚ�.} ���7���h�l�a���e�3��K7��O�f.]-�����R���^p{͉�F,A�B9z�6�:�v��g+f�-=�m#ڍ�n>�X��	{v��E���>q��5��6�%�*�Hl8w �x���9c>��?᲻���JJ���钋jY��S'�)z8aMOd ���_9$� �A�K*P�ç�%�0�C�j�k���g��7�l��Vx#>B�x�U2�E�)L!iA�WfFVV
"�i-��(J�+���}�P��][c�R�6z㪇���0
�XK�No�1��S��X��N�� �;�][@��2[[��f�+��л�Y��37�|�?,�k�ќ��F�9��T��fmTp���H5�8aDj*��ƛO�v��y�w	�'݊���5e{~�o���;+�r�؍xҿ<�����$R-�����5\��&�b
�v#WftW��<��[p��n�ڦ2���
*/���#5�+��5�9�+\B�B-�W{������G�*��Uw���I�?���I��s`����1l��`����0��$C?��G��Fz�1�����!�o��(���6����o�?s���������d~y��N���_�i�V�uI�T+ۇ����Z�$��F[��IHJn���߰�G��
W��b4.0z�9C�(1��!zFY�.�E���S��J�vsuS�FS���X��el�o��۳b�$z9��%dI	�\{�h��a��/�f
r��7j� �a=�Di��{rR��x|�PB�uɉ�4gb�ѹua����фM��i���&�]�u�C/��%l���9�u�]�Qͅ#{��+w�%Eb��q�y�Z���֒r��F@V�́�ZX�?B$&A����);b�q�wOшo �Җ��wp=4�&�H�;� "�J�x,[��W>]1���^��9Z
q�4�#��*���/<�xz-�lk�X͠�d�m-"�D2U~egg�Diޟ��O�"A�V�u��$p��1G"ɏ��e�jlI������%�/�8	�v@#��Q��d3�
!R��&�Է{��U1�`0���c+ў��ؿ~��������k��`�:S��Z�Z?���cX^�u��~�C�V-����Oo�3�'Oi{F�y�%,�ьϥq�
�f�Ťi�Z�t>E��Ǻ���e���k\V ��|&Jz�Z����~px�A�t8��j�X��B_U�;dO"�HU	�B��"�#��K��8ǖD)_���m�+�����D�2�f3�q^[��+�r�<`8*��(�1U��!�N��rQ�K���O8��[e)������A��
�2әg��7IŲJ`,Kn.M �A2�K�+gQ��/u��=�����k#��,���>3lH
��*��Al�;P~���2�\퇡��rcL�Qƍ���&����$G:*x �վ�G�FF޽�kb>H���"�#����Z��l�L��Zϝ��/�,� ~���MV^5;G�\.�(�|��:��L��]k1WL� a#]�]E	;1���r3G�Rр�HN���6�)�H�)j�Z{�@S)�E���0�O`����R��}ɤ#h�tKTC�1y�ܼ����͟�#�3�*��=4Q;�= �N� ����7L�<S2�ng�`c�3�o���d|;�&=��Y��ʶB��a��b<bq�Kx�ۯ/���
b�	�P�w��_4�H��ף���zގf�Kŭ��7�L?�� *;��bo8)�ai�Ծ,��W�4d�;�^H�`\zlj���J;d!vR%x'�H�9x۬Ko	q�}�:�l��T^�x�Rlx�=ҕ+�C}�g�����6;G!��z#����s�!gERB	̪�O������mO��4�`h����P������8Qwuuh��	a%)�Ņ���|��������e#ł�ԫ0}_���^��T�l8�� !"��� |�v��/����0��e�`����vo6ǣ@Yvj%tf�"�6,TJ�P?8rބ�p2]`VE���s�uQ�O���\0<vƥB\�K��'��u���?� 7��&~orf�����;�O����(�*W
![�V8�U�1#�WrJ�~E��᭏.��#VO'u��J����94�}��:J��m�Pp�v�����l� y���ҍs=�c�(��>&�֦�}j4]5Ƚ��[�(��.��.�ڗp�B2$���hLgm�Q�;����5��Y���?R����E�i��@�{+��t
�E�՜PJ~,�*!��W��[g�E�y�[>T.>&'\�5]���Q���iS�`c��(���|D���9��Ѻ���	�����^�����R��w,H�Ԣ �7h���7#���N]��:�@Zo�����ږv�4G��b5`}n^���Á(�P�M��$��ϵS�@!�bV� ��𱥄)'���"4�:H%�غ�Յ���3�]FNX	o���G���ŭU�n�6"�ď���-'| a���N��bV4%a�^���k荰q8��#���,;G�⑀Z�8'FӍ!��4�P&C�O��V��(FD4h������T5��/X.Q���1N��|��\���7�����0Ho�U��"�D�2�Y��2���3@"�リ�!���|���-�����S������,W9B�.f) dяf���Kmb�lw�V��Q:���+0��f&��%�~?�(p�E���g
=�WC�+�m��Y��c�<�[?����������t�[2�n��u:
 }��m�b�>��S��oG��E��!��4�wPΌ'YUޝx
[=DW~��Q���z�Q�EV�%�x1tgaoͳ�:�ef�����8�TL<�f�jB�*"�H#Eg�k�5T�"U��E���ud����ut�͊V�\�:�۳���i���t���{�1)�q��[^�4�#�"��U�vq��s8C'*O���E���H�-%�d_ә�+�Kب�!���:A��e�.�h:�u5Ooٮ�˫�?�n�&Jzr'T��^�ں�ڛ�9�l�P:���.f��aȜJ��"�{�*�7):F��G�XڂҌ���SaM��*��+��+�3ݏ�,!�.��~����	��qF6*Bg�A��G�2X���h�~Y5������F�Jpi�u��%S��'
���`nE��4�$���q z In��'�i�Q�*V�������IM?�|���V�c(8��s� ��ݧ����:���
 8>F��X��d�Y�|��#�����]�ڒ����a��P���ч�ͣy��[��;0
R�_!�iS�ˢy��)\,� Q��cX'����*d�l�ǌge�w�1�z���Z��������e�ܾ(�ي���e��x;�#\BVX����Y}}����������8W>��[�|4M���4T�"���_c��kc hw�.��c���HAJ��o CL�M`�	2d����D��*'ڡ.�h,^�E	���Z�*�Z���m�U:�S���S���5��e�A�W�VΧ+R��f����0������"�'��lB50�fQIQu����$��f�c� ��[�&����g��E9m�867	�pA
Z^<�S9>�j�|я�g`�sE�j�0�Ҷ�cL���$U&�F)����@��q"5���b{��"4f�!�?r�T����|����~B��������ö��͖.P��{�M�����F�[��:�8�"�;�}� {���%8�2q�&�����+s�4K�7,��^*�BuXL՘v�F}#����]�h���N���^r@�'1��Jgp)�O6B(�f�@�Ҁ���] �S̡fwOE2�.Ҝy�cW��Y�@���7�u�$eum��k�� �5�~�����/)�2��SH0�Dhy>t"zF��M�p�56��0�D��w���E(2�<�|�4�G��$PH�4�,H����
�û�!E	ֲj�(����6��*�7D{��
��IIC�&��C�����&�}&^,,1B[�J؆�����C��Y�����"9Ju;5��]|e"���� �����}�֢�B4�f���z�bf� 	Y�4
JV�f+"!>!�w-���fb�t��A�<pB��s �ug�����xOZ=��E���b��1 �mA�C:�޾5cfOZ]�s�������*dQ��5��v���ʈ$��/X2���ȗ$��qoF8����Y(�oI��J��y�Y|��(*nô�7�+c#iK�R�[�6�Ϋ+N�}��Y�V��^K���Oj5v.��X�MI�q���$��;�NV�k;h�n4�L��7����2儍��ٯ,��ߛ��DDP�XxyN��]�6W�l�@-6 \&��H~�J;�5A4�\��m	�hw��%����l��c�{&��3��)�D�wkvv؍����^�$�0���1"W�3y�1��W�dDy9P�S!�x#�/t�8���}1ZL��aF��_ڲ����������ڨ�D�̘��,:�_����v��(�ƛ�U��.p
���Y^.I�{���e�y}�UyS���!Z��5�U&j|��ݚp���ԀK7$>!6E�y|)K놎�Ȼ.�d���賠<kW�[��t+��UfI[m5�8	���Ƨ��3+0�7��f�%�3p��z���1dPx�	��y��|s/F���2e"�+���	��'�?7q�r ���\R��O����r��&����Y�7�6�u��ۺ�z%���=kX�!v)��ծ��u�f������E��.�n�����[�(���M�������0����v=��qqI�)���SÔq�m5���$B⤾S��bI�g������[������Ђ��j"m�?���dp���}�^����m��M�{�#�8���i��#]-98#]�q�E��%ad��7�g�.O#�Ԝ���_���<��*��׿N:j����t�������.����wH��$�9��"AU4���y?�-(f���������'5�V2@��ʣ�,�s&���|���f�Qֈ��T�c=��� �7 ��b�E�̨9���9�Դ��$i��2{����IB��+��	%a��.��I��릇��%��|�>��+9 j>0$a0�!/_O��	�	�i���ec��0P�cѨ=B��H��+�ql	d����Z�l�Eb�h������y%t���	�A8��8���6�ޑ\C�O����y{�h�� Σ�ӥ�?ꑶ�7#���C�L���;�\Xg �� ��(� �~#��'|�H�h�ao�1B�yĥ5aG�|j�ɓ{~abF� T��Y��4��D߻ �������=A\��f3�>��%䍒+��9�ݦt��1�<y��	~G'Qە1̆�bH��g��Jčpj�s �t �j��Ů\��8�H ~mR ��26��w^�	2�si�#A�a�p"����{4KԪ��V�5
攏�H��5δ�0��l�>�4e�~�\�[]��T�&%\�"_�O�v,�6�A�1���}����Oe�g�'�h�%�+���[��զ���R1��ɉ�5�:7Ы�M�ʬ�Ƽ�&��&І�(	l���H�\{%�9�4]K�B2X��
X����@nR"�uj2r��`8��,�wҤٟ��$�+����5� ���4o�~')7��d�У'��1�0/8�$�}֠��ʳ`C�?�,���~��{S�Կ�M)b�W�3��۵�y�!)����3�ԇ�Z�ȯY;Ɇ�b�1�/XP�
��#	,Z���Xt� �V��'�:��G]��i��bE���$D���KX�	���)����Ѩ��d��0����M�(�V�@����IH?}�6�)*�=��)���z�-����#��{K��fO�>�N�N��R���������P`��=��
wxTRm�T���Ov2�P<�&�����R􏼈�"�+��Z���-�Q����[-n�A4�`>$�x���R4;��?���?�:��E�u̽��o5C��m�IϦyܯ� |qq
L�`G�]J��Z:�%�3��`�����F#�"�V ��A�7q�W�G�'A6Z� �:KT?�B�L�5w��]g�N��%>\͇8��I����l�P�S/`}�iִN��y��Ny�Z�a�YWAY]��,5�k��� �k,C��C�@�r�
��s��*�jM�vɮ����e����緭����d~+e*���eG7ܭ�fA_yi%7�w�D��1��V�(j�	�����dõ�%��֊��T� ����v^�u_�dAiH�nʟ�ȷZ2f:����Un�X%����R`E����c�b`��f߁*�[�m�6��	C^ak�1��`���w̕hi?k,C��OJ_s�3�O��N ��<�V�4up��5�	ؿ�`�l���e��eh��n<Z��ͣ��g��(�loD�� �c��IX���z2?4��㝃����ﵞ�1=��j����5M	y�T,]1K���ܱ�wo�����������s���� ���jsQ��M~HB��4t@���	U9�=��@eA��O��ո^u1J?,p#i�e�y9�X��O�P<�y:Á�W��.,�gXz��b)�͠g�O��8�p�c��rTr���YPA��1�]%Ы�.�s��
l�6ǆx��7h�D*J��__ˏ�%�p����Pg�A���7��2RJa ��m��0��&"W��e#t�f,ǣZJ��^���0��@���$b��3�16�`k�K�ٝ�+Wh��QQ���ԉUR��JF�
�%�_�����w����K
�ǣ�^��	�z��+ַ�ɘ4��}�>��C-���r�ئ�X���t�f ���LF�t�m>��&�����4�H�۱��i?�ߎw�H}�)x0�%9'���0ns��,n������-�5�'YJ'�����s�*�_��.���J���S�Gu�H�����I���W�|%���Lf�ڣ3�"�h� �����>�H���g�$� f������u���P3@r4hVy�M�M)��2���0d���3Q�?�\�6=&����8B��(]ȗ�q48Dn�ہ�2K�wWY�0��]�4�C������h�.��9�w���[I�/����9�%���o�����K�t��Y[�`��y~8J�η{��MJuN���x���1�x2�g�<�dWc��$�F6���_cvi��6j|��t���m�m����E������'��J��Ӽᴐ��H�_b�����3nn"]Q�0錄{��,�쨪��0������|���ƭ�MMd����yF���Ө}3�ou ��<x�A���[Dv�x�s�ȭI$	��{�ȥ�'�e!ە�7d�lgSj4��bᒾh�����u��q۴�v.�̆��.
�N(�֭����<�v���&v�KۚA��L'�����[h�x��x�'ۧ�X.���0LL��uD���� DY�����Z�>��N��g���,�ܶ�E���Ǽ�:���ྉ���y,iu���z&N�9ߋ!�d��꧒��g$���l�}�R�9*�?Y/����}��o�#��5b���ߠ�������v���}%!���%���D�\�^|mKz }��
44�Hy3��ҋ{�!v�/�R���4����j�"�Q`ѣ��t�FTF��>)"�:&>�����i%�;���M�J�j��'I�e���0����:�sBR�D��Z�+(�(x�
R:�8�,�%��'TOE:Ъ�%ޫ�?]"A��*��F��kZ����9��I��Ш}�T�)������uH&F�蹎
~(���6z�ō�S={��v�W�)*�d�׻"��FtD�c�eCf�t����F�yn�$��/=Đ�
x�g��U���'��ފi��q��C�_*[�-5x�g�����9ſuk&�����b�q�0؞����(�����n j4�d{���g�F�XR�W�{vcB)�q����1��Rvڦ;������gP�˂H�@&�+��A�+�&D�bȁ�֞��!m�!a�W�߳9��K��C:�&�p�ϱ��&Z���u�ZN4��^�Yw��Gy�ҝX�(�tu]ׅo:���������s��5F|nI(d�b�k�\=��Լ)Y����Zv�La���{�,W�<ի[�E��XO�x��5�(�L�_u��-�9�7;*�><��<z@]#8�\��a�ql�ٸ�K���U®0CS�9u`�OjO�YR���'����p������Ԝ�/�?w+�u �*(6ҹt�J�6���;����&�k�O�hZ�a�ߟ-n��tp��[�TG���T�*�3���:�j�J�v찚�?1Vx����Zz��'@g��Ɖ��X@;�U� }`s
5�����߇}������u�]�߼��sڠ�1Zk�8?|�>Z�žcqF����3�� 4Ar{�K��?غ��V��2Յ{�?�o���q�n�]�]��#��:#˵�i�O�q e���E��V<�W��L
�3V�%n�]��n&���#�A���ƥ���X�@u�K��i$���?�A��n��J�OS���ɽ�[ ��V�i�z����3�&�zӁ�;�h}���e��i���^�t��Tľ)���:-.�S��/��e���=3��>������\VBDZo񈷷��	l�I+�Zh��z��	H� ft�dJN��Y0����-�-}�����K���g3%�!������k�͔�h�
M~t4ث���j��0,�R��')	�	�M��x������R�reN�����'e������MD�h��J���(�)J%��	r'ʮ yF���H��;�Tf�-���%D�$��>h��4*SExe�)V��t�ε����>	߮﫲h|UCf8�����\'�[y|�8+���D��2W��U����j�&<X�O���S0�W ���`��)�� ��'����\\
ˢ7K�i)=�<r��F{��h(�()�w8������K(躑�4[��hѡ��HK雜Rgp����S���i����zs���N�:#H�;5�0[����;	)���^Lj�i���ѼԠ�n�^G:���]~5�e\2{όUq͹,(���`k@������+E��J8����u�C�f4�(=!��oc��<��ԣ�%'W�r=�#-ߋϏ��"$�}�oa4%3�xh�×D�(W��s(����Z��H�AY�u�^��߰ld2jP��JTz���3`^e{� e��FU�����}�&Ҥ�x����
�d�^@t��p�_ҵ�V�L6ҍ��]n�Xī7�{4\�%@�2��Vd&H�3X�ޛ�C݌9�|������o�G��t�/aF���ݩl�Ȫ���3��NQK����eʀY�i���I��rWH�s�/U4o��鳬o{���i�錁k;���У�OW�/�_4�����c����5�y�`��~�T����k�E�����p�&��8?�J���Y@�`�) �W�ѝ�M)#@�q�cd�ݽ��1]:�%z���hF\�vr,�����n&/
='o�'��|{��";�'c�E��"�Y*�d=E���}�Z��(=��C��i���-!2�9�/�i�a�\h�aJ0y㧪���R�1aQTȒ�1>|)�����!9M��O$�G�$X�
B>���\���j�ny����#��5�}�7r�W�yy���X>���-���6Xk��bR�0�i
@z����pkn9ǪW���;�c�*�a�ɈT�������p�i��9�P{��8��:�f��O�͘��׫�:B{j}LO&�w;О\�b'�;�<�cj�N��ºSug[��E5ƽC�+CpJ�m<���o�����d	v�}�/m� �b=��/Kϔ���]6K����о�s�]|�Me�̽�����6{��(u{YR[YܬQ��ڵ�s�Z�qkK��A�{	��]O_��#�OM� �G�\���b���Q�xB�
�ǢuH��:��ZFs�#0���H�"^V�׵o)���J�4�Z�/��{ uIѺ�h�4b������%+>���iۡқ�����}߻�C�ӘAWJ�tJ�;�OU+�	�p���Ys''�1i
yxg�}�Ʋ& �/Ѧ�b2X��R^�o�`.�0K� J�ウ��S �_����� ��t�����e�@F����2��q|�;�6 ��?>t���7Uf�����JYw.
�)����}v*����6�9���C�*G2��.I��ɐ����������n�(��I�SL��٩d]��O�/�����������Ch�r{YT��\���T9����-o<*��b�������g��#���C��t��+�3[�Q�N�N������I�Z�5@���(�ُ����*&`+o����N��%9�K|�B������r��<b�?_	��Vs�#�����IIPپG�����d��CqΓ�/�N�TCxQ0�#'�G�&��x|��Z���
������Ɂ6+EsŖ������A?�V>Yj�	��ܗ�%g�?�꼐i�_�\_�W��K�UL���.�)�d"¾8�4?�<͛�>U~jiĚPW�:!����ٔ\/�J�8Oc��n�:х�EI�ms鵲~}�]���<����cG:����r��h��t����6+��X��ΰ�wi���n:�d�]!~�Qxp���(T��V5���H��7Q�!����#��@�KW"/ �~�g�x�!��fp�I�G �D� �:��Y�p;!�7	�nM��D���܍_@K�*���8n8�7�y�*�18��g��s)�i���`��S5\�T:��|�`����Ue��O��<D�[�'Y�c�ח�:��g4+/��M��Q�ը�L6�,Y:x�U#\~�_@�_Q�����zF����EK�;֭G��Oz�L����8u��qn��S�=R�y���n��O|	�L��oR�vX@�~KphU�|M-�+4r�u~$ߋc��\/��F�~�RG�;���F�+ӯ�i��Jx��|��JE���&�6�s�V��ީ�̄~���<R�ڷƭEc����Ѓ�_�j	���}*��?8��$;%h�)o9�ΰN�f.�(�h�
d(�8[�����n�y�rgXz�������o2�m&�m���׋b8K��O���OÊo枈�W�M���P��j�ڟ��]^r�Ȅ&�,+�[DH�j���e'�"s���J�lA��#w(L����^NꗠVjLv��#zO�asѧ���.H8������Y�1{N&^�9c�
�T
7��f��$@����n�1s�m��%Q�v�N�9T���3��؉z8ᜮ��)6��2�#g�l
B�(�������0x��#)w�D�{����|�m�ν������`�<�j"�����<�eEtC:�~5�L{�P�v�Y�w3�dMR�m�-XTZ"!��޶�bf��$��*��q�i�����i���("+VZDLz��<��|��օ���s����g���(*q>�@�^āq?�qr3��Ym��[�CDS׀�:�{Υ�#��b�Z���;=^/�@�������p|�>��������H;�ģoy��m���6�w�>v.5.�?����)��`��,�X���$�Qb^�	k�A��ҹ_����(V��8D�������)�kx������Y�v��ҟ�m�6@�坠mk�A����9�Fo7��M���?�\�/�$Փ���){	�ɛ��-��*�?�����`���e4���n�AK ~�6��@#�P����V��3�n��g�kƈF�8#?��*�T��&Y����2����m���n1���T���`CLF���dd)��ء�^u/�>���	9�^�w��0�*�B��h��׶���qg�~��cgGLexDsxB䥤W����n�jz��SG4ac���OU��i �jB�@4Tk�[�ԓP�ut�)l�_)�K��W���H9^�9v]��H����;Vo�܋TܛR֦�,{x����pw}�$�suRD>�o��2��){gF�r�����/ BL�j?-���.f��gԺ}�� {Bd�Ż� ���2�(�!�q~D�@��}��É�i����e��У"N�p����3��h�^�9�(.�K�-���sG
�yRk��њ��Y���{:�J�9�hVt8��Zt�2[��5lrrh8��m�}�Y�xcg���)_Ē��] M7[���e�\8��~�`�L5
�ogv��U���<�Ӣ�z��}%�- ,wo%Ȼ�F��f�U[���_��7T���ʍ�r��8xƭoK�=!#~��r%�%=����M"/�W�X��ZJ�����0�A�M���>4���6�����,3_��^���pM:�2�,;zS�{��1S+ .��n��%���p�7$Mli�f�+o� �3B�e?<�r� L��]�?r`��J l���`+'??���,�UO�w�*�3Y�?�VEG���� ����,'
���� �pV�bx�6��E0�o��&�w
��z��#R��N{ 3}RCGguy��*l.(p6��P��H�P^G�fz/¢j��c�)���9j�4хW�Ѽ�x=����A]~��������U��t>NǽD.y���$Laa�\��y��k���3PH�ؒ���X%hA�C��(#܆=n��.�"v� ڮ+�y~���t�{���i�tt
��/��g�rH`�-U����l@�ٞA�G���R9~�����;L���T�e������3���<1�"��k�U�1�z�>5�%X�s��ϕE%��aC��޲���$
|�úE'7�UN�'ulo9��:���0L!ǿ����� i������.�հ��Q�'C{����U�e���Ag�K�ŉM�(�1;�)A|�<m����Ed�@٣�C6������j!���
/��WL�I��U»���%�����>B'���\��Br�^�uD��R�Py��".4�g=4�(��Gl.��ӯW!g>�)A"�b��C�,�Qя��M�fΐ;E���q�������F�ciL8p̴^^��&���4�&4�2�	=�Vvqh�@/-QvE��Ulʀ�� 3Ƶ��$�S�(�6-����l����@_�"��1zR��w��8����	����z��hR#K�BE���v*�0*�l�)�X}q�cWp���~�0pв�^�ϐ��足�/e���[�\�b��G��b�,\N&0W,��Mm|2�R�`cɱi�n*�TA��:z�'6[⫑p���?��ř��x�[�u�x�`d��V��G73��-@�/;�����/Ï������=Odj�U�nc�P�
8ub�|�5e�-�d%�[��f���]:.+ϱ��$L@}��cS�R�3 ��L��yɔX! ����󟎼�����&���Zo�5����9�GC��`�b�Pp^vs��7OG�ٳz������qD�Q)V�� 	���
7��x>���$��ń��GW~K���,V�7WhZ-sͽ$(���xЁ����1.�i���d�+��c*_ѡ��'��Ү�Q����Lh�_�������@�Kbk�����d��m��q�w�U�7A�� �EƔ�K�|�X �Mq=�"�EK��k���h�|o��Z�����[���&���O���lg�a�x|�'kq�Qz�}\��9(�����kCİt&��S��m4�c��+�'� �P1��66�F_9������mc���I�@ ϰ:��0S���ṙy�\3�,-�S��~�&yIj�n���B���C��"�ts�vR�b�[׍�Yņ]��k��8l����46}���i� R�������w�s�����������`.z>�UD�� �Oc��H:��ٹ����K�t��̨Ѩ�{*�d�%5/��U��������PN?UUj_��'��� ��G8mS��tëN����i�ߋ}����98N�ł�:�w�k=�P�x 8@��s�/����|Y$�_���f����~>��į/��µ츈�|��&���N�{W-(	>і2�.�0,�܍;��s� �r���b�	 g�f~��t`ɓE�I�ý:� +dǢ��?��+���΢-��$��C#�ރ�	9lڕ0�_�%�n�� � ����/h��$wl�R��Y����	�V�լ\��h����w�xH�R�yPLV�ǫ�Ok��d���#F�Z��;R���TK�(��6E$/>�m�T��@�I`�}�M��:�|��Xz=�Coz�8=�>�zK�B{׳�I���Ŵs��Q ��U鋽��]���Θ�N��RԼ"PK�ņ�d���&FQY���=���K����Oz�I�݃�E����*�.��Ւ8�,�
A�V	�'�%������1��YHL�s8�VY�H���7�����?�J=K�A��n�_�G�céh�Э*V�8W#X*E6�%���e(���Y�U:>�Ę��*L���ג��^޶|p����m%j}m���*]"��$ؙr7���g�딟���w�pk�ۚ~������z��)������R�_;P��Fչo\ޑ���6nԣx�[ؗ��5���������z��h���`x��1tw�����Ϛ��:X�Mc�R�ן�}(�ʆ{C�3���p���������۩�����lu@��J˽�<I�����o��������a���I� ����^�+�,�� hY�P{j�,�F����.{��w��D}�cLCD5yƸG�=wb#�ӽ<p{��+n��Uɐ�R�����>CP�@`A"݈f�u��&Z����j�1��m�*`vo��~={�!�N�{�,����'4��b�ְ1b�����i���a�ih0n+ �4/�{��aԏ���6�w�CQ��,˱�N���ۉ3&~r� ��T��j��/>reWM
��Y��3���A�'~!�jpO�E{M�WU�X7fmPƏ�Tdg�=�'ֶݲ�Y�-�m,��'���;���%=7���uG2n�3�o癗{̩𖈊�3��*-�aꢗf����T/="Ϣy���x`�V�XiE���9@�j�qw���%����w1\�!5����~���0�k<����<�_�#D�`���޹���I
#���eޭ$uQ'
!��Y����%������H�*9�Te��V͕GŭjӒ���Ϳ܋���,33��e�.$-��|I皱i�@�����"X�Z,i
i���	�i����f<G3zS�h.
PA��T���'�(8��������JXl46�����[{-B
)<��QF���t��>M���+�2,6�^�g_O
~����P%�΁ډ��B��P*�:L"��pf����8�x$?j��B�g��>�R,<�w�Vgl�����$�b͑*�ਾ���S�Ӽ���VW��?�ģ�1�0e��U6��%���w��}G�����=m���aP LG+>�^���2H�n�4�v\�?v+���:���9V���&'��߽���+��@�JY�Q��$���A�{`u�7�^��8�������'�?�y9��?#$<�f9ʁ���r���H�:�@�,O�;�!��S�qӓ�r�L*��^�y��g��E�Ʌ> l�����f]��?[~���Zf�r�6P^Z���6���i�DRM���	�(��T�h?��!��e�w7���l�\�m�'[�j�|�u�9,鵈����W@��L; a-L����P��<����(��[�pL�\i�J�4�V��$X��!�Lއq�Q8;Y*+���[�d(k?�l�����c�m���{P��
�}��@��\@��@��D�lw����H ��<�A���1�F�Z��XE�O|�L�jz��΋S�E3rà�׃��k
�]�}�3*�x�CJ��8W���f8]����r�x�jPv�Ofi�`��-�e5-������w:�)ȗ��e���թ��(���G"�^c�|2\�Qa�X���G}4!�2S���|��ٝ�
��`
)Ȁs^���aV���ܐF7[�H����a�M�F��ȹ,K)e,
��n��m���#��z(�1��`���1`�YߵH�j��φm��trU���rHV)`�
�?�c�8�lBmĒ�骦�.�+��	�-�XZ�>[j�w���������w��7�΃�����g"c���Q��6�$�?2qs�r4B�%�L~C�r"F|��]XRa�0<�ğ-�&A=ye�J;��V2u�e4S��D��|��>�)���s�ס��Bq��7���
�Dn��-��� �e˪��\箲+�|��Ƒ�W&�?���~�G@���Q.Ҷ�m;KU�;��a��9��N4�Du����j�kܫcnt}�%�}���:LL��-4PW�ٙ���b�7r+|��,hK�ڕ�_���N;���c��e�G1�Lu���	]���[2�z�*�՘?e��IM�Y� zQZ1���'�+!D�
?D:(9�T�OdVsX�i�6m-=�&����ڎ��@@���P���|���T0��S9]��x5Sq0O�&��C;�Cǭf��I)
�z<�e]��w�@HCU6�kcN���`�TK��=>JaE�{\3�"*O����D��o������?�R���``�>�s2I�	�tdr��7?�g�)�D5)���W74䯥��X��͓���ö c�d0Y�3�R�䥥��cg$��J	.�0#|ǒA#�:Y4��{�;ε�6��\#]s6���Ɔ�4����$�6@җ�a�I��=���#�Edd����.\zG��0h��Qع}�,v��C�P�:�_�=�A犿�-�>�{��``8MH�Sx?�?)�^��{��О�0�0�q�Y��I�ݭ0w߽�ӛ��;F�p),CbW/1sm�'p �{<�a�i�
��'���s��MM U.�Nt���)�"�'O�q_%���E�R��LD'�i�e��
<w{��T���=R^8��`�_L��-W�*ԟ�Ѯ�vΦֈ��Kī-4����t�e5��BI3��]jGn���t�8��/!��m4�NE����~������%�W=.����@o��%m$������ T����M��Z3MS�r��.����t;��1e'ɎT�G��F�}Z~L_�q�5c�y:�������,��V����o���5�*���N޹�x<b-��Q����\[]��$�����T�[�w�,�����\6bn���V���p�L��,�\�NZ=a�Vo)�?�e^kU~X���'|IN�$92�ը�J��ڻ�#�E���Z��,^�j��2M�F`gos�?��K����V����t��.$W�%K[�?�FG�#(!��e�?r���x�����K�Ӳy��f��u�K�|���ў2�nuׂ����$���T�������I����e��)-2���{{)�[��9��uQ�Ǿ�j
Xg�1S1��&|.g������E�za�K�i��:P+|�W�5�f��@=R\�c�nF]�kۢc���o����a�܏��P�D�sգ��"��MԺ���P^�O�orI�E��;��4��үR��]O�f��z�'�r�=+�g��)�<�X�aRBl��ת�Ufe=A!��~4v0-�<�!��E�/k�H��<E�_WkE:�Svl�T,ِ<�>�h_u���O�y*����ʒAeGE?��(�hՏd���#��{�=��t���"�T���a�zW��Uw��S�������9���3�U���I�O)Ad�Ly���R�u!rS����>�����k�-+�}��?�o���1��������򃅪�L��� ��~L@g+�?Ӄb!�=`MhGw%Y�uE˵Px�*�nx��e"p�>�w���1�S��?%6�g4V�T	����:���"�M2��d0*�R+�>���v�w�`��8��-��쪎�&	�������v:�:IjUZne��w^����Y�3 �YQ���_v$tK�"U�(Lt7�6��J���7���^u/%_��j��V����ɴ,'��]�.�<���%���6��5\=���]�H�Å['�D�k��(Lx����6�?uPҤS؁a�A�L����1�ږi|"��7,<jc���h�+��/Ӿ��Y@G��~�fD���*<��!O�ݥ����31#vaW�
~c��wώ��*4��I�'s0W,�8�o��E�v˧E�`��'��8o]9ێu���WL
�#�5����w��xm��E��VQ)���C5d���^��*9�=8��`n��q/@/xLe?浱M��S�L4"g�}�jQE���P+��$;M��u����V��.��D�4�o:aE�d�	yO�G���Zuy����?�����g�Řc�X?/<��R:p�	��!�&��/Cv�������U�D�z�;���lb�K����01w&��������aR0�KiE�{y嶈㩶(?���MW_�~shӴص���91��N��}X(*�>y�,}��������7A�YE�GmU<�q���^I%�mj?�w)�ƆXu�xI�S\�(n�ڱ^ ��Z������Ӥ,?��tD{_�X]2��}�FM�=�	'��u��ɕ$�kj�QNZc�\\��2җ���3n�W� H>�85�)��i��f�d����r\b��5��#����/�?Ӗ9z��������oS��[s�K�ޤ=={9�d>�*����xL�K�P��(���HqϚ*S�:�Jx�(��kk�Z���s���-�+-U��~U7���͵��_}�$7��,w��v7Y�������q��"�G�e~�ӷ ��h����=�z=��eQ��,�LQ���(� #WY�pw :������V4�$��M�Y����ړZ��J
�,�z0~���Y&�v ��EѨ�71tM�g�#�-�)MA`�/�4\K��i������e!e��F^���{�. �"L	V�RT����v(�(n�Em�5�����Y���j��ެ%��+p�*m�c�Ը!� ]UFS�N���h ���<�0���W��)�ih��7Z�4W���T�o�e��� �1�B������x�<�� eH���׍��ϫ��#�z���9�`�7V=W*�U�|��Mǲ���m5�5Q$B���$5M]�CK������ �@�ee��{`鱝�4�;���q`��e��V�Y%��>����l�O0 *�����V��Φh�m�<�+7w��b��{�0��+��/�����.�t�/�����dD��k�6��?.�I���Rf�δT��c�2�T�M���$.���W��ph�s�<�����UPo�*KT�!M�%0���zu<��'\��XM#��0F0�	�G������\̣�Z�P�4r��+$LV}>�̩Ⴈ�=�e��[,ٶk \I�0��H�b�{w"Aﰳ	���ל����@%��ˎ��pM����3</���E��;��=�3����F�d"X3?��.��r�f�4����Y��mlJ,�}bQ팭xY+����˼�����@-�WQ�����j���ʡ���-h�Q'���e��B:��a��b���z�c����.�DS��0#�h�K�� 5��wZ��_7t���Ȳ��3���?��o�gI�H���,<����a��W�<jVs�)5?���N�5лo�[�C�b�y�5���r�R-XV��_��%���^ 0����wDx謣����Rҋ,�y�F�II� /��j}���7����PZ �U�Bط��
1����X�e�u���v�=��6�� ��}~� �-! ����9�C�,�,��dǧ��M��^cŃ[)��~K�i0Ț5��m���.錖����5MB�VP�~��i�l�s����s������ϿW�ͽ���ŷQ�3�y�}����=�����	?��ezq�d�~rF�.�xS�Zϣ�� �"���Q#.Rq��v(�Ǜ��UJ�0�f�S
X?Š�va���	�^�Heʟ}��`�3щ�I��'9_���Jn=]~���@:ѧ8^;�G�:[��t�Dos�&uF�K>��zv��9>�y���_7&��{o��	C|�f��g����������P��cg~��w|��/���0ky�R'�{���,!��ʺ�	d�WZ6��WQ�:����]h*�9�{*�!�K7)K��ݣIl�^_,�t��eh!4R�e� ?��X�Z ݟ�e�^^1��ɕ��8e
X�/F��_֦�"C�Wn��&ԑ����^�v��t��t���2�M��"o^-�w1p"b�~�ԹB|&� [�Yro�2����in�7����]�#H�-��5͍Z�\�ŦOޤ{�ə������R�j�p�s��@Iȅ9$oRm�몈�Nh���'#⍵��6�oD�Hy���Q��uTGD[rXM��7˹7�f�����`�f��@���s��e":NF��ZgK��)��,w��x64˄�]�@��P�����O�fՓ�`���r�Z�!��W]�� ��%������uH�Tu��4�ڍ�����v��"x���x6��%̧���7����n)pˏ����������ӓA^sh�eN����'kKL��n�n����n+��9y*Q�S���K�M�Ց��:� B��K
5�TѴf�P��"��!�V�d�\�H�_�\�Tyn*�-Z?_�)��h-��g�+��h�-v���-R�踽�����~=1�.N�N�x�jo�u��a�.�6f�?�Qg�~`�پj��\x��˭!��+�=��*�4x�4uw���E��_�+�M�����_"eQ����JJ�\����j:�1�r�F
��
tk6g�ÒT�f=��#�kH	QN����1!b%t�G�Q����"l�5=[	�e��1֗�_�~��.��
o�&�;����sꔖ���qQ:ky���d������*~#��&���H���y�\��R�J0h�H8	�AB���"(b������݆/��Iq�C��aL��4��� �|���l� ��<0w�����4O#�5�٘ w�F�}:K9q��ez8�'��'_1Q���Eg8rX��h6�����v0h]�q�*](K@���
)�)[���ϾnK.�rIB�d��tFρ�����S!'d$F��Z;/�K!6�ƒ"TT�`<Rs���#��O$s� }�~,����v�?'<��d��}���!�$�O��Ŝ)�J���ʣ�$�lSU����4:$��̓����5o��,�1N51�ՀL�D�Y�{P~;/3�/ş̀�w_�-���o���Q�(#Z�6��槫\⮨��큭%�F854sR�����S�M�]6�@%X�@d�,][B΄��ꔾ� ��E�sZ|]�LBu���@�%�As����u/_'V�7e�g]P_�IJWd��
}<1u�ɴr�Fǆ�T)O��2l�m�����Wi)��R�(���*q�=����k|��^Ԣ����
�����u<�ن\�'
uC$�ڣ	�Cb!��`Ƒ�;Δw8���ݶ\'�P#�$�7Pn�u=�A��V%�U?���bI&�Ͻ�ɿ�:F	L����*��Q>�b!-M�;d��M�l��IO^����������'U�.�Qq��Nq���:X�;����;Q�Ƕ�4�#"1�R>KX�׏e���M��������@S2"Y트D:vz��/��<"�Zm�F-����7jQ��ﰚ�^�C�O
�@���cc�IPX��a�!'m�A-��F�]��D�_f�_��ͥs9&����Ĭ��(�)��X�!����|j�W��fΚ)��1zS�h��|�;=s̒stv��}���h3Eu^���f�8bc�-�6����d��dF�S�3Lj	�l���ޏf�R�͋�c�/��!;K��@޹��L5��
�����u]��
�bo:��J$�o��8u����+��Tw��&&U�^/
ܲ��_u"�	Y��ݭ��C+�Ws���	���
� ]R{�.�H��oLj1��Ɖ%P����A>��`@�h�$��C��Uᣢ��Ǆ��{��(5�k"+�4	^��bFx�9
�U���ҸaV�Р^ch�
%�8{ĺz	��T���i�<����m���n�Y�+T̀����9Eĳ�"$��],��&����l�P����Ř�YN����f�]�Z*$� x�kz@MPv;���B�gI��z����B��Hf=��9��5����]-{L8X�b}_�,a��8n���^9N�\���ˠ���{���K�~�{��r~\I! ]b1���[� ˤ	�] ��X���F*��ªg�ͤ-�#��O�ɧ~WA���z�ڪo���z�d��^���k��
I�|�'^;O�\�m������| ���Yz!N���Og5�L&Q��ՙ^�+mf�J����qЪ�2��q���Y?�9un�>�u�M>��o	�t[^L�l�!���݋��tZ�8`����L5����R�>{&�Ƿj������~Gc�-u��QP�.�]]PP$h��%Ά1n���R3H�}���cB�/������
�~���/��y��%Z�]�G��[���\�ܭ�bW"JA?+1�����Y~(�r7OC�6�R��$���[�wQ��\9CA<�����>=r|�P(�:�fc��Hwۈ�K'RN.��S<�=}nD�/��`�t���s>5�����&�1�RLML�͑b͟�<G�,�?(���yqQ(a`T��ԙ����А3#("@dJ����I�`��]B/G���6Ռ3�Ҳ�9��L*�ޮ��QN{O�"<����@X��k�6�v������0�?�;(�:��o�H}
f�i���JM}�pR�u�}تRuI;���$�g�O^AL�?�.~��������D4]��Yz�ߠj��6��l�e�Ϛ��q�@�[I�"��뚆������3r���݀4��$���&�W���)\�=���bF\�Ky<�g?��^���)���0/�;iF��j �\cr��1�U��}{ÆRTŐ�n����4W}��iK���1�<�I�b2C�\\�eo��w}A�" h�G-Қd{���(���ڲ��O���	���/M~#�T��x�ez��l�d�V���j�l�n��Yw�%icf��W.ڊ�����:ol�n��mK���I
���8��9dF!Y	�#�K{�MpXf\i-A^�"vNвY8�}�z��'A��wcȜQ^�MIKQK2�/v��jK���^;A�w�G˽3�����*����:v.�2Ax��a��.{wiy-LE��	�Т7�Z�����X� �P��S1r�89n��T`a�PM�:�����ٛ�Nߵ������X
�șV3�b
�g��0�v��.�n���w@]k��	c��^�-M�X!���ۗEH9�$G�qfϰm�y�,��>@ �R^��x�,"��^h2���8�k����7d�Y�2EAz��~o_)�b�O�����H�U{W��CDb�U_�%!�m@��D'|&�r|�J�[��Ιg(ˤPV �"<�'�6����~��P��=��Mz�!�M)��iq�p
�>��Vwَy���N�"~Rm�/M�sBx7��X���,I[d�'զ�'q�q��n���GvMuղ M���7�%�A`�r�c������8;�:�ke�@���L|sr��-t!��r�ȏ[��
�­�0�d�8�G)��	�cǎR8͊_HLZeu�7Ve}O�J0]kY��a}AM�dn�a6Vδ�Ġ�;�ye���v-���k!+j>
"Z�mu*�/�9rfJ¢pw�=Ž>@�I�x�Ih����ﴀ閇�`q4��'z2�֬v���H�4#�.K�n���Ke�J���`B��ҋ�{�<�R��e���:�����F�gh�����t�♒��r�" ���6��ޕs��y����^
_Ȍ`�#�c��ܟ���1	�;=o8<9p�4|'^W,�Aa��x�P 
�K�b5��#��e\aQc�-2m����+�s��;d]|���8.���0-M+�&�kDuN*X��4��1x+^��{1pfO��Al�D�9����~�����)����Fl�{�!L/��lm`�3��b��[�(����Q%ah��`W#���럅��Ұ'������m�_ՏO��'�2�Ť�6J�R'F�6`Fz�|�<�
�c�o��!g�K�r�Ļr�+7�~�	P�FnM澶&;}�}���Pe�a"�����)8jt+��:�,���W���{�d�p�9ҋ�AXI�v�81
�?��Qk{�~������I�}�#�'�����ﮦf�eu���qa/\�� ����E��Sc<*�4�f� �/��m���nl�ڲx0͉�z� ��DX�Iv�gd�ǣT�6]I[b%k��,��i��a��q������lm�%��V�k�<�1I�����+�� �D�;�X�HD7˖$��F�g�B?̷_�4�Gڿ���I�#�=��n�*�	����zo��q���,Pӆ��un�Hf��^[����328��X��1�f������n߽����������8S��%���C Sݳf�yl�8�`�A���i7ˠ�x��A�Bse/�n�?F�J�=�OH��䤚f
�0�M��Pc�埡i��K���,�~3m��.�)�힍lo=b�,���ϒ�L+^�]���"�@Ht^2��2��Di<@ �ˈ��t��S����4��&��^s�x�y7�=��5:�c64���~��Ǆ�x��L�q�m����\Ͽ+u�G�:��<�`+����0n��;~��
%�	�z	m6��Ȏ��C�XP�_�I�C�m�u%[ؒ�q���X�%��*jJD�P;���0H{۝B\���eRǾ�X�� zC���� ,��Ң;�=�ړ�Yt֯QR�3�..~U���o%���@���e��R�g��8�٫�ȗ�o�~��la(�29]֕��8�*��!�;21�����H�K��)����ߡ��hqw�K�Z7�+!�2�֓��|1e87�~z/�Ԛ���g�=N8
���ՠ���
�N#����D��ͼw/���f(G:��e��lN9|��(�-�|bO:�N�;	"°��������J�/��q�(�[�9��(�bD�9�^k�ft���B*�]Y��~���:}�OQ�!���_�fƧ]�nR�TZd-�� r������^Ҹ���)lF��A5���/%���e9���m���r��Ʊ�4|mc7�i��{�_�#a���R$Ab�"�J�s�֔�yݘ��D�N�Ny��[b��^����}0�75g@7f�//��<7�>�g�}�:���~�\k�n��t~d��~���h��.�x��e����G�u���2�F�j��`�O�������~cP_��:9�#=�V��Q�wy�B�n4���O�h<�R�٦���ͤ�Ʒ��q�x�#+j����4��"�GJX�sP}Eb��z0�хN�;��'�O���VPM�x�%I���&�U��L�*��ل�-�7
m�q��6��68�Z
�wd��XLQE�3P:�_8�]�Pg��z�
�b�9f	a���clz���nk�����N~�0;M+[�F���Yyk��fvo���g`�?���Z%&tI�۠'��5�أ���xcF��=&=�|��20����h/~O�`H�k�It�B~w�Յ���{��[�,��5���z
{+��=�灱
X�s�,1pN�a��� �Bh�ZԔm")��c8�a�N�V��X�
��q+/�h�M[�������2�BiI���b�?,��k��<��T�����&��5�O���hmQ-�Q����./p���C��O"��l)I��u��c��r���A�|�Z�Z$��[��*�����Ի���)��^������CF{u���@bS��9�����r�#2��uŨ ���_=��e,��]Z����Dr-��?�������Pr(�BN���mAu]l�k,D�����z�p�D�.!�DK�����ޛ�@l�� �S9�F���	;��v�5�9QCj��՚�����gw�avm�ͭ���@ϑ�g�}
��@$���19	IːN��{!���/��0��M/���"��7�(��������ݶ;�H��,Q����#�S��� <̓�,�P�Q2�o*�@�+��}�𺶥ۈ����py���r3��ŗ�h���}!�WHLN2�
�3�y�}ĎC���\բ��	7����(�������럠	;D`i��� �p�&=�7����q��LNmq�m߇��~^]uɎ�ٿ�E�P����N��8D��y'uS0�p����/�IQ��`/�z\{��V)�b�fM�>�C�g�s��Qq.|��e�P��[��JB��Bk����49�֦1n��d�
C��}8�$S	��r��[$�t3���9����s#"�*,%�Yk��D7��R�p���u��`�
{�JdC�4��֬��P\�d�:�o�b����z�W����ņ�Tx�P	v���G�E~�x��s{\  ��y�#���-,����NN���͜�U��Y������Nn��(�7�J�u=�b@��c+v�li��c�Y��Z�x�`u
�yY�0U��5�"/������2���Ͼ���=l��ﴳ��I�+�kO&M�3eY�%�[�r�M�����Zd���a���)�i�'v6��}y7�31�r��&�ޡ�{p�o�|����5Ѧ_#a+̐�@�ɯ%и!M>N��w�� �a�X��:;NC��݌��o#wGG�z2�S���I���Xt�.( ���~[���곹�{E�ЅL$����,K�7X�����X�;P��G6�*Vt�������j!=�s�%� �4�C1�L���[n��Ǵ��cj����ԟH�CtV�!�S�G h��,Z*�l؏p�G�NKH��E	.��U�0EE7�=jJl8L^�踶q��<W8O�p�l�ҝF +�������.�q�-��7TZ��<�~
=�S�S��a$PZ���h6�B����᧧G@����|ބA�h�M���"�T�����fJ�`5b�ե[g#o��e����e���[5�!��ҍhMlpRw��i)�~��PA��)�`
6N�͉Z[?���؏ǚ�8�uZ~���ߤh��wR���X��H�����dk&�i�a��.�Й()��t(���eM{� �2~0�i8?hbG��5����4���O3G�V��Z�x[
��0}'_H�g�̓�q撌����f�0$�פ8 ~mË���|�Xn1�L��68����I.�R���f���jʼ�n;���|ΡҏJ��?��&�BXqW6ab ɕ�ԔhNKV�wɈ9�;�#7�Zߺ����y�{����~~�����DG	\�P�Uʒ�f�����p-|2V�/�lf��u*;5n4O�g����@H̚y�e#%���\�'����Q���oE�vS` (���PX��IKRi	I�R��0�?c�����&�x��m]�u6�x�1�y�GD�SZ��R�9BV{��V�ͧ������v�l=��{0�����pؗ	@bY��ͲR&��-O�3(ґ�.��+��L�K�d[Zɟ�Pa �c7����ڥ �������W��b�*�x���.$����W�ʷv�cՀ9��U��`t�B2B�#��-���{.�a�ʺWa��E�x#����X�=�C�_oL�7U�LRvGײ#T�W�$58ىd�>x*$�ؘoH��F(U�^�/���;a(?j�0�5~��C�w���;��/n�Y�!�� ����F�����#��l�?��D�1e��pZ~B�5lr���d�)X���	�jC;I&�5%[��pj��a����/%��רs��8�M��Z�6ј}^k��d��qv�o�����,�#��uTv%JAb�c$o�ץ�x�eU����p��*"Ql�� �(��RX-���el�(,���<��2��E��[�0����T�]}��vR�]�k*���D��3�h�����E����,�$wޟ�����^/h�i�
P&ţ�8��}=���|ȋ�㞮R��Z�l�����Z�H�Fs*��]�E���a�/�܍�I��kkqk���U�6/UtO�xZ���������E�{B��H�.=���iCЩ���n���:0y��W�0��-�
(��d�I�g,:}�8��6�2{�6� �G�	;i%�{e���z�T/ޥ^ț���8t��W��+�4,eo�\X'��<-����E ��,��yW��͍��!.d��E}��{)�V)-��;�"�q!��@�TC�Jvt<�*կ���� 6&���ưS$HJ��2��!;;��ݛ�hT���}g/�V%������ �@yy( ah�H��]��_0���
|�L	�OK�Mƈy&ؕ$42��>4�6�HJ)ROd�kyk�G��}���5�� 9,;e����)��+�cp��b�h��,+;}ճ$��v�PZ�Nm^>�`��y�m�;�'`N��}n7G�W��|��c�����f-O}�4�ӄf�D6n��*PV�&�uפ�H��L!ٛ�n��ٚG0�'F�	j�`S�H�+�����T<W��E�4'�4GlW�}3���y�T��{��p�BQ�1�{IU��"ɂc1� ��s�C��q�z��PN��k�����s$���W5«%�g�oB����Wx'H�2�D���O�!/�^Re��yL*{K2"^�v��԰���Ҙا���~�Rb"Hs�3e�%|�N�^��s
��6��,�q�\�i��0��ʡЇH;��?0�k�nH95�ǄӟM�w��T�u�(�w�?��(a�O��D���<@߫M��}P��bz
�V�fD�a�����I��o]*�pB
�z`ޥ|�<���\���e�o����Ym�s.o!��CD\s�BV�r�q���I�;��G���Ƕ{+h]j�ޘ�&(�%�A�#���h4ڎ@j+����o-@�"�d�-�u��N�-�F�;�GB��������N}�S|ʂ����}��u��S�Cj;ȣ�W�������wƽw�W\1�q����M�4N�Z�!3"��f�&w�d���6rz�\��g4�
�rGHC�(BD} �(����]F��,&�Ն�f��r��	U�W�"P�������D�@0�\��<��T��S�,_��cRB�V�`Q�!����?�@a��Br�������J����*�.	�d�aK4������ Oo+1yR���X�	%`���6=+��w �$��#�N�w��ލ���LL2��5��X|"x�]�C�"�x̫�������2܏�/��z`5F ��E�
A%n��М�>u�
"+�v�a�H`l�BOWb����5��$6䱷�U��0��n���g��nl�H��1h�#X�^6�g���N��C�D��̍��zA�46�?+K�{�:�.bޡ6j��lӳ�{��|��m�9�q]��_��*)c}s }5���M�>�9n��V���� �u�M�J�B��[0�ߐ��48&c�4�`���3��M�Tk�O��s@�L��pm:�K��~���OM��.��.�$����dH�]�H��$�O�|ɗ~��<�g���у���{dR:&3�S.�V�-�@ �K���{_��/���N1,���S�J(���b0����0=�1Bh����P�P���`3� ��݃Kk�*�ֆ���*�-y,Հ4{.Je��2����PȎ<�Ɓ�
��� �}�� �6�C�i\�~"���Jk�*����h/i���W�$����%fؽ�[�Hc&�0�%T�DѾ��.��]P�оf2]��i���Mo�h<
d��}��P;	��A�r�;E��hk@E>�;d�2y��`��_X
���вZ���"e>	!�E�E�-'=�Lw2e9�>q��-�M^��8i��'��:T��|�
9X��Q3�"�nt�c��-'�_Sz�G�3�oJq�o5
��L|P�
()P�e��3�����w;�����p�gٜ"9��|Ig���Ӝj8�����wO���U�?M���ڬ��6F6:�C&�}\Jl�l-�H���I�j�k�NJ���rۓ�gRemd�o�h�pXc2h�@p���o}�,t��4�'YDm�m���%�.q��k��B��H���G���Y����CV������f��IX��8�Q}B�	*O SsU��g������Y�ҺX�	!DƋ�F�(+� �_'��H�<�Ih�����I�2.R����x|������~.X����G!����g���ꔡ�Y�]mO���2z���<�)AF	�RcD�8i�>��`������tef�~���L���R"��40���2پ
��P)b5�����;�+�lC�Ȓ�/ْr�a�
���/�qȖȒ��{�M H-$�y)�vI>�ה���r��c���)OZ�+��2kaΛ">�/T��c-����)��A�XV^�H�)�)8BU��[��A��'�E�Ƙ/�4/�X�L7�L�������P��w�l@[n�Y�T c���n�E� ���>�%�u�DԻЂ)��ʒ�8�aVH�|uB��������w���l�ڶ���j�	�MY�����A�p�jf�U��/�w�1`U��Ҟ���%l�;�1'��܍�(Ph4Ő��Oy��1����S�����]-1��o����R��cb�3��K�iFW�n�?+�����{f,k=��
������Ǔ̮�ю�J���@���uG_����� X(''�������Z�^��Sb�=���l|Ê�>���/��O|�%����S�8�I�$����<���=��@�8��H����NH��L�3�4�*��r֕J���Ń�u�e�;/��S��|�<_y���^6�'�Q6�8O�v �����W��;:��&�]%i�s�m3TY�6���Qt�w@�/��˯�؜o����B����ܖyH^.�a�S�n5�S�N ��#bqeqP�8F��P��DN�z�E�Փ�ѶHI�U�3��^�r��i���q��#0Ɋ����+|�^�#�Z���=�ʟ0y��0���@�%k8cz�����(o�i�Eƕ�#Y��i)y�j�����ۑ�N��j�ռP2,J���a�&.V�5�n"0�d�Ϣ��ciTU�Ƅ�C���G?Ti%�=5�~���@�|˟�*cg�3 �V���@��}fB)	��8ƌ� &�����Uߑ�˺�3�A.�������U#���Uݯ��/��g�pE@��Ch�ڛ��>��2����,��O����e�����҉�o?�t~|N���z��{/���~�*����O�v�\9� ��5l1p����En�eI�b�Z��N�.ܶ��î:��6��w'
��˧���R���s����k87MZB$��T;4���ϭEo�j����Ю�;6�}}�/0�oh�o�|C8�1w�cc�TG��}C�k�R�ؘ ����v'��K�zr[�_�}x+[��R���O&����h^_2R�q�8 F5��t/���#+o��&��ip���A�Ay q�ǜ����;gC!E����ˉ�+�[:���/Bm�U��3��ICbh�	����\���*TM~�������p>���F+���Ip�\���*�?��c3�! ��Cmk�ϓ̫�9�<Y3���y���oZSi�boƝ9E�h����sx]�,`�.���qX�|�kױG'Y�L7��A�T�0?�X2���̕/��7�vb��S�O�#��
<ެ�&	�ӟ���QH��@��7�O1F�FY��[k*�M���0FK[����H��K�폵Q�̋���ߕ#Z��D�m�r��#|��EFLֽ���)�fP7��X��i_5�������m���#W�]��(�n���#|^�J�[6��z�����Ӌ=��K�;�* ,��mG�8SH�a�;��Gu�µ|�xg��Kͤ���A��~��ls�.�}t���I��5�;���W�$���P�cs�ӂ)>��Ƶd3C�����Q+�:���'�ui=ˬ���A��ǂ쌌��ȁ�'���Ĳ����4�^�Mkq��.���ͨVC���8�x�G)=��X��U�c���e��y"\������n�qriU���4�=&�\�����s؟��Dr�:�#7-ΰy��Q��@J�^w}lQD��>�V̺܄��[��u�l�`�m�ad,�67<�4��ŜHM(O�A����T�`/�p�Mӱ�m�0�%���Ne��)�fTH?�2��#V�<V�J�)���=&�8P�^H���O�.A�m�z�d����	_�J���y.�aɈ"v9�E�d��4�u�+���j(V��K\�=S3�>����ι���	��D�:=��d/�e�X���DӦl����zW3�qǯȎ��M�%Lg���Z4S螖�Xt��>�ޅ[1�#/�o�$a�ף/?�����Q�b�=cW�t�����
M��=��0�bM��յ
~�r��>���d-ғy�i��ug��V_���k�%�L&3w��x9�o����%*Q�b,���{�Ee�*nco���w$��t ��g�re���E���k�s_��=Qi��J%'���&�լw{�Ը�u!��]{�%����$>�8������%Կ�ӥ��lh4������d�G�}�Ń4�N�ն����F̇��}�Rȇ�F	)��a��2%'�#�S��	g�Pj�;&����rw�,��$�H��P�T��;��z6ۜ��7���}j1r}�<O}���K��"�mv�Hv� B UxTq���k*!�'��^�d�[J}ﰳ3�J�lXp�.�J���^(.P���w��l�64��ڥ�v$=��j��$E/50���%��Vg��$j"K	��}o^�R�O�q^`��+U�)��>b,BY�
p�4< ��t_enc���B,<]gF-O+0���y�3�������"��%�6��g�a���t��t��n��u��k����{C�|m���Q+����ʺP���Yi����\��j!7P
�����!~�# �����mۅ�y{z�C_��$Ѭ�S�;�8|�!k�T|L��Y��c¥0u���(�e��)�_�ɺ��_���U���2%bu*��1S���Bw�R���T�"KH��u��H����,���
���h�(v��w0b�$�([v���d�̖�G�"�+&ѫN:e]�����]�\�.j�W�wQjCG���I��IUƻ���[�p�A�}n۳�����ڙ��6޻��0d`�R�Y2R�&�Xo�'���jE����Z��6w�1�(��/Sy�W��|3S�p�Z���l�b���^jsoXoUA �9�A������p� c4�2�|�+��_��JN&U�JL|�x��LM�i�}N��o��$��z 
*bP���#P�S[��j���r��e�?}I��_ԙ�C� �g�(7l�b��ih��4BL��Q���������l�K��n��2�s)W�G��L�[bx���`s;g��w����,UZ, �,0-ص^j��^`l��g�Z�#�g+���jCMML�Ǿt|hDM��jih���IJ�za,?�����:W��5V��P����Ǳ�l�(r�Q�W�0{;��Ϋ4�v�L<�V
��T�U38򦇟��rdm0O�i4仠A��UVػY�t�Q),R3��04��{�W^g[K�Q��Y=�B2���H�xB� ���5����gh�R&����CN�~��3��`�|O��`t:�#r��D���u.�Z��@��n��H�����m��s���>���QK$��>�Y�h��i��O�a'M҃��Tv������T�W�w�*F'/Y5-x���`#3�L�'oTG�	�Ѻ��=J;��� ��~Й'M}�a��X��}�pۥ����Z��v`�Sn����F���ў� 5(�f����hP�a�H8�4��`g�Yn��5G �3͂��^�P�Y�Wm���6� ����A��ڧ��ƀ�X��9��̛����i�t������>�e&*kmؿ�Y_��Y$���]��S���Λ�k"��aH�H��cO�-�����f�<��Ƅ2�G��Hv'�s�ҍ|������ޕ�\��	��>0��q���}6>w��"ž�tCKZLo�����B���P�瀢k�Eg_F&ǅ����d�a=�?#�jlϖ���?���M��T���poP�����Oc$.(6�e��Y�C�Ҷ%. nJF#�?�C��P�\�J2v�OOM$�4��_2�T���=�>�(	\�q\�C���~����$�-@��%��tMO^��;~��ڤwR�eyꞱ�*ɝ$����ȼ��*�cԿ��;�ݗ!������r=i,��{��	�	�k:�)(�F������ �v���'�ß�Zl�ϼz)���Ĉ9E�I�O�:w�w��ЩB8(�� Ʈ�����쳧ҩt�8JymML�!�	,'Ha_�u��pI��.Ƌ�]���4TY;����)4�D,����R�����a�^�L�``������ ���/%Q���Ӕ 
s܃�����]by�"'�!���/ce��u��m��8�\o^CM� �0o���-�B}�|��Fn�2�,�3Ղqer9y��yiFN%�Z���j��VW{��'�v�Ώ���sQ��D�j��3+Ґ��u�!�mK����]l�(���]�uu_[N|{O����N���]�(V��2�U���C��࢒��GG�,n��	�����h�
y]���F�A���X�l��2 £_ٔ���������ӆ���ӡ��Q֣�͜�覂31�p�n��>ƮV��@1[B�A4@��k��bEJֵ�1glc<z��(���QWdtnsߢ������Rb��{��ξ4B�)wE��ù�w�Ɗ��i�O�S3�'N`���/o~i}��)&ؐ�������M��xц��a��7E�I��ʤ[�g�
�����('8��_��DqD�������!���b<���cL�J�ږ`U��W�'��o�Z�h8�
��=c��/>�iVӑ�j�` ���?�i�W�X�ht�'t^k&��od�R�aĒ��;:��/�t_�d�J�<Xx�D찉�&MD�D˅�EY��D���^�2AG6]��9�ݘC� �MZ'��:2�i�s�2�C u�N��L�^�m~7 $��a!f�5��އ��9p�)��;bݛ��*g�脗Kf�*e�ͫ҅W�H_q�
Èwj��=1JS�Z3϶T^�@&�a�ă~����:��K�d�c��q����V�/��z�(a'���۷^:	��T;��iN��������D��3uM����M�GM�@3�)�'�ہ��C~���#�Z'D�ؼl�=�Ѩ�	��DR�1��%���Ǉ���hֳN����l��%�	�W�k�����mZ-��rǶ���)�hT ��������m�e����J�	z����oy'21>��wS��u�V�ma��w����s�W0w��aF�Ư�e�ΫҞ9-�<a�`�=*�u]ه }�7XA�6U�|K��?�Pe�����ݓ�0GS�F�X�0���}�2�k�-�(=#�\���UB�é�H��L������.Fml��d�>�s
tg�Ie�<j���G�N��ւ�J�2r�d|?g�>_ך4�9�+.�o�S����GMB�1��h��wp���<fa�-�9N���$����~�(�r�ZP�>8k�W��4:���ˊf0V�"�X��#)�4�Bd�ݘ�Kf����べ!���QnT�&�>��^@�ܺu�l��/*|�ٚ���W}��S{���P�n�����ש�2�v�b��ۛ���Y�/N���2��AL2�p6[��!0�P�&C�!���c�I�9�%e���A���q����o(t��ܰ�j*lKƑ`�!L<�$��"�,���׏�,����,�WI�N�שּׁZ���ϴ`܆MRh���^ϳ���x�	�/�Ά�$@*�k�"�v��:���|(��tm�9����Cn��K���j�PT��$�2��2ѮG���k�)�P�jAG�c�R-�9��:ổ�6r|�Sl��$Д��k%2|�a!�Ϛ%��X�������❥��.� @��e1LF �C��v�
p�NC��=�jf�V!�j�@�؂��k��#fCz;jF/Ko�~�q�M�Ss>:�w��c�~
�#=QC�fE4+U/W�������gX�
�����n�D|��e7y�Q5���{Y4��F��M�%��{q�@q�ҁɢ�[3���1�'��kq=U���ځ.
3
�-s�AƴߜR�	�ؐ�RVP,o�?�Y)�ק��3
p���`�6��Zr�9� ��4�#�	_�ต���\��S@pZ�ʅ�)'T���2�<L�܁��-�y
(��[���*b,CU�:s�/�c���Y7;A
ϯ����|n���� L�ӄPa7��k|/ǶȎ�oO?�P��Lp��yT�[��D���|V%A5�1�F��H�������|;G�3�r�eEa+�!��æ����@"0i�i6p��فt6�Wڣ'���b�L|��c>�ڗ�̎#S�mb���#�p�G��m�˕��s4���@��侩�\��K��X�DJW�܉�D�-�%����6d��o;��y%��/���sܲ"�\q4k��(��k�52ꮬ��	��s"\P�&�kc�r���h%�UNt���Q��O�b�iٺq_��$�g��Q�n�r���0 &F�7�gY�>j8�@�o%��	��pZ�������ą�\C�ba��*�0� �LS\���q�*��C겚h��%��� p�����kz���/��ӦY}�&ש��C~{+Z�[O��)�;���/�0f��Sxm���fz���v��	��
���ފ�u�ڹ#/�nI�3��ɔCFo*�e6��
rj�$Ҽ������_aPO@�pΰ�����i?��~U�x�B�xq�٥�1ﮅF5�^{6�]�տş٘�YKV+��<���_ J&z4����5c��|N�`ƒ��Ɠ�'7]s�83�@����OZo]��>�>MТ��'���kI��*ҥ�����$����԰�Cs�O��C=��C�3V.#� ��a�h�y�~ !�U]I/��#Xjܭ���Ij�:�0jȀ'T�V�J��
R<5���O3=^�Sv驖�&�	a��k��M��ۙ�Kĸ)~A٥�im���nܟCЈ����I��"9��	A��s��e�y�o��L\CN��j��!�F��|�.¦|�
��Q$��f.�c)qPGe nP`H����/Dh��Q�&�Ei��d��7�r��eE"|���*����7x7�Ty�&@��� ��OB7[I�pA��~1[�̌��/@S���L �괿34L���ɾ��#L�#�=��\�~����xE�- ��0^�6�z�,�w�n���`���ڌ�*A�?���}��ƞ�+��oXM u)��?סC���Ȯ�ò+N,�F�9���I���%MS��0fA����:����A���zj��f�6E������Z˃�Ët�m%�h�SU��h6[)�WYob��'1��]^B���@���O�:�&�w:_��.ѯm�0'{��
��m��z�s��n��Ň���Ӭu�#~M������{o�Tb���E��ä;[���#[}q8X<���Q�h�}]�P�i=�x�g�<�!2s�'�	���7�ߴ��s�ѻ�}��OV�M��j�{�GFq��w^�>j���U/9U��ޱ�%a�]��02�
h�I�߀���"�r��@%��a��V��PBR.4��w`�B%ЙՆ�&��V�"vAݲ�(ƞ�\V�,���=�5������O�l��-~���J�;6l`�(��x�)j�I]�-�91�>��C�vF�4� g4}�^4#i�*��żiZ�9��gI��e���y'����ǉ��13X�����E"vZ?��W*z4����R��(�ű,o��sSܶ��D}I���@��Te��j$���$�nkl��{!lb�l��㳿��r��
�~������#�����~{��NS.�@*��df��k%�Z�<�jS�*h=�$g�.&$ߊ��li��~0w{F����%��z�B?�f>e~U�A��<Բp�*�v�c�dd����I-�Q�[�n�;<���ؙ�g�`�~h���K9ܪ@��fN$tbyښ(-c(`@�v)H_K�� b��?shZہ�Q^F���RO���� � �W$w����}R�����LF��lrCK�<w	a�e�2ű1K��Q�
,Gt��;��Ovp��QRU^·hX�õ=��鼏�-��A����2f���vM�Vl�cE�2�Å��xh�������� �����_�	�v�����B��ѥ�������C����g-#�ص{$��o
2��3��>U�YIQf�j�RB-��R���@e40���3Q��yʰ$Y���~�ɮl��Cu�.�i�Oũ�궝�uP�]٬ݮ0ňD~�t�3�������L�/,'gLx�E����4BP�i��8�B�-k7l��Ci�c�@����ȸ���xw�mEA]�\\�-:�b-�I� K�V�7�pƂcP����4�s�b|�]���q����宏����4;#���&�R�[Λ�hNЙx��B�F�F��WU��-�kT:u<���M����y�lD���^./?Awю�;eX�yw�[&m��
�R?&�l�6�cV��r����jMu�}�-���,'clw��"t^8�Cx�o:˸��Q��;Q����u>��T6�c0x�vjU������[Z���8�ɽ��ŏ��cr9�D]3;,��&
@�D�x�l#���PeA\����]M\�h���2�Ֆ Kza/ЏE^��[ݜ�Nem=������Q�tc;w��̱����l�wF�\�z��:Uc~w��_�H)�|��1Ϝ�����W!�%��:�e�v?֟�����r9Og��,SS�*��ƕ�98H���f[)m�[/��e�������i�ޑ}t�I�dh.�����͆�S�_#zE!���tL�K��?0�X�y�������H8Բ�$�����i)�i�L/A��gS9�!?�:�4E��|�,Y����wpň%��1�n<|��.<�z :��v����2a����FK&��d� ��j*��Vp*
J�'y�]ݨ��������2C��w��������={w_N>�C����,�d���'@��𙋰H)0�۹c�	�G�Y�#\�g�R�M��ht��%��HW�)�)����v�H+.d�``��q��0�6���j�:_���3�<ޮ,\�_�U$��&�����t�Tq.��<������ܤ'��_�a�#��e�]��W_j/�����&u
����7��+��p��k/#�m ����v��1�� ��>ٖ�jZ�Yω��Li�]Zfuν
Ұ�L��W��B	���/t�m�&�W�Sw�p�өY�7� �z��_��E�uah�fB9�$��0� fX�'�qz��_�a�M�`Aυ�_V�D�O�l!���q��n�`j�i��y��KBru"�_�x��^��B�������!˚�w?Xj��
�_3�Z���=�R�����$PIK�GV��Hɴ:�y��v��q��''~�$a���~�����c!q2F�U'뾍�?3�T���Py2��?c��A�6�I�<�i��_6���ӊ��>?�z{<x/�y��5����{k���r�N.T�G{I�6�гAc2�n^����ܧ.M�Z�7�@�n$3�>v���+8�/�1]w����j���s��5VpPᦺ�t�l����h�?�D�Ϸ����d�%���D �}�d6R���J�Hi�c�����d��" �ݟ��c}�
�B{�+~��%���J��260)�6���7��6bV�tw�a;\��-���a74'֟=������t�fE�C㬜��˂ �F�.���/�icr3����X��Jk*LG�?Ue.)�����p#����G����	���~�-��� �ekK��ǂ�7{�����H������~�x��yO����O�V������n�5�K73���Hi�+L�c׍��(JOCG톹���I��;�e�ծk3���>OS��7�q�-,��gg�/���&q��3fH�t�D�vo�V�*�{��.-��wA	�ю���)Q�Y޲����l���Lf�Q�s:�������4�޵5�Ծ%�r��
���>ŘV��wx|	�u[���J�t)�'n�l�=��сwh�6��&EMݞٰ��q|��&����*�6���Fް����!�GMV�2��,��d<��D��yN�Y�@����Ko��s�q@n p}��OV=�O&G�����<l���az�ȁ���PS�ǖ�~��s<&�I�x֊�"	�x.�B�i�A��n+� a���E깉Xǐ�;^g	S��㾤��-~���V&d� 0#C�=��_�S=\P'�m�f�և��8j��>��3�Lռ��aN���I�<�yԕ!�ʝ2_|��'�c�GT���:�� M�B�����(�7��'�MOH���ڢ�����;�~�2~쾶�Q{�m��F.�����-��X|sD8XI��^|��@�1��w������(�5�b#*7��e	*_�LԒ�D%M���`�T0����4"���m��݂k�޶U¿��Tʯ)B�� �2ӯ��9��w9�N2�!V���Wy�
2MJ�ҁ�-�I��)Y��LM��G9��cCRy-�fR�C���o�G��n��;'N�~��35�c�|C���4�fZ���	�R������J#�Zm��� �� ��Z�L4��b֨�/�����+�q����ٽgM��[�SQ��B��)L��߃^jA�g*��.9��(�WNYř�R���t�at��p����N�kQ���y��m�D�!��yJm�		nCi�.�f�a�E�5�,�]��������H���N苂d���`�;T��af�%k�_%4�D�����F�����`�|6_z2WtY`� Rl��!��g3�-{�A��u1mg�ƭ�LX�?"L~,�C�5�F̮7|��:_���bHi��8B.��hf�|Q?���f��'��Z��\'�ZY���K"��Ȇ���D�z�n����On����XЪ�*�����5�'vle �F�[Y����"����w��ny�5>:w�"� �(�+�T��x4�����v���w@�F�Q5�"��������=O<s��Icq�Åޖɥ��k�XH<�B%��?@�┢ŧ��2D�{�pV��3*�@��rJg|$	�okH�ʘ~��[e��1�ýb�r+��!j;<�nLho�GI�
`��i�����E����4��P
0�bσc8;����ͣ[͵ߢ�3��7��1!w��9��t
29�Y#C���}�ԇF���~i����D��hl��Fϋ1ه뇰 �6�Ԏ;���^�8��x�pr����I�>���ގp�m'c�Gc4��S��!��S�6���n��T�9�ȁQ�I�tx�(��0�jq�8"������L���64fw� �+ZA\�����~%�ŵ��T�q��-��~U����H��v�#���YҊS������SVtʍt����5Т�V��7 �u�3�0��~*�;�D��#5�OK_���v�]8LS1��o�O���8b��,��Hg1d�Y�%���������C�t*�l��/�J�Cm�}	��M	��\|ؗ�����ľT���(�US3�JaV� H`՞cz�XDl1`�@G���T)N�!l^g�y�hL	G��~�a����唗z�e�Yﳀ�S������:Nt&4mi!�T
�ʚ�p������5�͒���#МJ7
V���<��Uf
O�g�t�/���aǧ�!��=��M�.��%�&m�b�	���'o�Ez=�\�O�䀃k]%�r�ӯ�%��n��H�M`�pO���F�2�2��%������L*�m�GSk�ܮm5TK`� ,�������; {���}e��yƏ�J�ՇXu_}����c�<�0`����ٍ����ɒ�g�7J��`�x��4�Q��~C�`�n�R�S.��L���<�!Y���dG1~۴P�`r\���4�.�H.³D&�Q�k�l�l+�J�`� ��%B��FŒ���K5�L��8�>|ʭ
u0�l�Y"�y����J^�s	�=V�Cyvk��w�u������ŀ�3���H��.�7��� �j��zHv�u�}����h��0�,����:ǿ�Ǚ��Vp�M��<m�a�$'�hM�3p�)��q���nR����@���Ot^�Q����Y[�m���`��nc�+z����@N�֘*�������7�=3g����ztl���bG<w�g���0�ci�[�f�ԛFrDx�P�e�}h��
)�4��ytq��v�.���[ʯ���T@�U�h�[�����V-��'�So=g�W���#/JlKtws����oL���j��k �P�ČUUU�ve���/1kͣ�ȷZ0W�^)첑z/��U�������cp�$��?�Z\�?�/�`��Ç��P����ϩ�{U������ۧL�n��`����K���6��X֩D)E��o/3}{R|e&_�X?ś�w?k���	i�,D��\
��/wyJ���^F�%O�P��ᒣ��(����y=��RxaT�-g����}
˲�vI�(�4G]DE� �9�z>|�7��hdΦƕģ�t�'鮯�$8�T��<Mv��y&�L�`.�,ye@9�# ��i�I��p_�(�혷�Wՠ���li%>�Ȉ\K_S��lEą����Vg=�S�rFO��~Tڌl��Z��s��oBX��߮/�,�j��e���rJ���Cq�����^wtn�,n��}�iy�+��N��io���B����#5GF���
���lW��^�U5�� �~JwI�U��;$��e���\����o�
I8`�:P��G����}�a��$���L�Kk��A�NǙ�}rA<���Wƌ��*���;:�JV�-��6`�Ok�#���e�H��4o3�v˙<�z�#���]j�AB�sL4&����u���D� u��f5��V]�5��G�֭ƽB�L�X��x����x�q!?�HhaЊl���^��j�7��Y��<���$���]N_��X�� ��"�*G$n��"'�="b�K������Ի@Xo��/������躔D�w�S�B�E�d�*���So�f���	Š��IGe������y���5��(xo�C9D�c��ǵ��΢�Zs[F�clH����jC���7����e^csaZkJyV:�$�u�I�AMOK�Z�1�m����	Cu�l8[�6u�`��Q��8�Zp}��7�(oPt��_�%f�C�OXCx��X���żU��Р%Q�m�,�F���=n�Z�w-�|5�����[��~���C5?��⺡nv�{�sz�e<�,(�*� ��y�Ġ�/�v���%g��ZkfA��� Z��z�.3*���"/��-[��0�|���
N����-a8��&sz�/�j&l�zoJsjfd���m�d��ɿS��M�Ԛ$(�����ꮤ��T[f�f`C&���%�F�e�P���({PY?qڄ~�������������n�ga:��Y�����
JÕs����$����,��2���F<�����l)�[Fz�M�7�S�>�FD��
��9Ӝ������@��<�b�t�QX�H�yqg�	�^"��ij,���gHo
�o�XOYk�`��6A���%DYr��&!Ŋ��J��åWl\r����1W�T��D�zlim��*�,$>�!ڸ��a�n�t�	rϿ25֏��4U����?A�-��F�E�~��S��?zN�������^�P u�b�n�$�.3���L�h4%�:m�2+��UQ��.Q�w�"�Z�hNuPLp��BI��i��]��4���S���N[ �/�<I�z��U<ĥ���.�7��,ٓ�g{	,{٥fn�L�/hz����Lr�^$�5�6�"ؾ��`��ʘ�Q�zz`�l�0��A(�� e��`��(֡�,�pG[ V)����D V
AHW�S,������<\��*`��5^�Z�.��V'�����u8���z����3���ݶ�	��J��k�8mOu苷BC�X�b�{��}��ɿ(���ZoH��u�̹��sK�J��R�l=�tm>]��������C����h/B�{c���Jd��M1k¶pVkq&����d�eY�r�IUV�"���[n��@���{�Д���Hu	��=09���_E�-�f���H�C�w�k� �c��+:� ��z�q���f �
��Lie��wg�{�'�au�q�'42[��{,�(�@RTr�e���{�K+a�if��_�-�']c�����*���c	e+h8���2Oӛ�Q�[��.Q@<�lx��zl����:k���5pCU�X�-�����W���K0�BbG��8��F5�f3j�k��9ʄf(o��l����|�}����u���<Y�����?��ǚ��k:������W\�á������6��Ho@QC��t3��;���aKc��2��
�yr�3{ȶ��;����B��Z�"��e�uǷ�Qe1 �R��+h~^��F�$м�kx�s7�-���yR���`�)��DU�L�����5	{�k�I cA��X~̣�Cn{����u��;�6��yt��$�]������"Dt$��g�L��	��Wp:��T�\��EC��z֮�z�A\������DP�QzA�AAr���h�Ɓ"f�4IΖx�9�m
�P�S�"��W�C��B�n�lf��	�i~\��_̓Ǝ�gG��+o����3G^�68L�'�֣,wA09��m*��H�o�����u�-~�)��X�o9T�š��,����l3��:x�ܝ1����od�
O�\K�$r���ǖ��֕�!5F��~a��$_b�6���^�>{�����h���xV���fB\��V���cD�Y����9R?׭���3���`hԺ�U�+U�}�f*�s"h�D=~�� W���+#�1�Y�Y,�b ���r��W���l�u��8!�M���6:t�P)�B*:���!|}7FǮ�e��p��<����u����}����p���O�8��r/Ѱhm\H0
;���;D������5؁*q��`Xr�����O,,��I2��D�e/�ْcM�ԟ ��p�����f�,�0N�M��]�Z�D��⊅��p,Qh����m`,֞�Xޣۻ֘�ꗨ��~�t��O�Y:R�A�i���S6���)ߺ =/�Zh&�G6N��@�v�%��׫ؘ,m�@�l�9X� 8:&@c�A/���A�ǁp�kb�6^����b@�<*��G�>�}��+�xvӲ�"RF����x�A~��'^h��V�)S�*��B@�6�{��
SHa3��
�6�RwL��o���)��^_���W�,Ϲr�2�R�ک�d��M�j�����&��)�.%��/�]��L�������D2�}c`�Rdy�2��m���T�"@V��|�>���,Zբ�2�����uu�]���c�_��+�����:��jK������'�	��2Ŷ�T�E�fs�鹀iPie�z��H�҆8�p��"L�+T�%�ԛ�y��&怍��j����)2Jy�"�G�L*��zY����d��ЏIo��(KAJя��oH�ʽ����*���ʒ</�?K�7	��q1�|�*�2fN�<f�Y�G���O͡�J8���h�`��Ku�Q#�aUʿ�񦗊�	���`�H���J�i����[P��7��/ޛF��iS	C�ƮLKP����\���aZ�<3�V���ǚx2�Y���ٕ����ණ2��$�F���/��X�Օl����]��IH��CO`����4RZ_koɢnܮL̍.��yu�3�KLQ���-���D�f��8&�r"oۺ�Ҹ_|@F���ܥ2Xh���~��ag��^O�Ri`��l���6�����Z��4���e�6�S@�y�U#��/^�����Q�A�:�3�S�t�h~.1�'m׵��;L��I,��Q��YH�.Ǿ�A;�g:҈ n��;�P�⫃�����ۥY�y.�5h�I`�_x6_�?����k��kg\\ ��ϸ��6��r�M��q�)R�Oˤ^�Շ�6���P�Gj/~Z��+�+�E�7�a���`�ڇ���� I	�Z�E_� ��@Y�O"��e@y(
?��Y��`�b(LJ6�И5�$^}��b�ִ��d�ʳn2,����+	"��]�B�Q�C|3��_�]+ ��8�C��ԉ�&��zH�}͎�� 7�#B�*+tӣUU<���q�,��u*��-�1@��*b;%�~q��rpJK��LN@��������1�HEW�JH/�B{1@r�n���fK���(%�f{Ԓ7H���r }?���oJ{:꜖�X�.i[�l�<,�\3k_��aVGy�Q��D��$;e�)�")�v���kOdΒ��ٻ�����.�"�[�����֓�/�̓�Kr��|������y�;Lnqu�N�[۱#5`t�RGHy������,1N3:&q�\=���~u>�����j�8,��3���>#����F>t]7�~�>\v����k��$7�r� �LA'�c����St��.�T�w�����3ւC*~GCA(�wu��^�ף�Z"
�0>f�[<����c�����;���	%%�e��߸5>����nֵ�Z	�#�=a�?��("�먪��v5�m������f�.���L49�N��D8& .�Cr��_]�m����@�����������f�l��	�g>X0�qg](/D�qԄ�f̨}챿w��ZcL�&tCR�`2'��Vl��-�E�Z|�5��,YU;�Y>x��y����E�O�E$ׁ}��0�hW�!�B��xj��V��h��v �=CP�+}��"4�yvRr�F�b���O-��-s�a>���=v����@�,[vN��j�n!2����9�#�E7��..,�>[|�H+u��I��n���4U�'�yn7~��y��8���[��\�Z2G�k~һ��Z��A'��=��d8p�el��;��l�j��&��M�b��;+��s۩����<giݜ2`VWM+4���BG�a4�Sv!k�{3ZU@�_���Y��ᵩ���O�!���MfF��1���r��73�g3~T�u�(3ĸ�K��9y̬�C�ǃh	��q�y�bF��<E����]���Ϯ1C3?����@I���r��4�f.k�G�#%U��Q�@Ϡ�7d�{���9F��?�\�M�,�"�A܏�,��2z	��!d��BKJY"�6eu��!d67���c&�欅�<���2�]+��Ԃ�ȉ��>�q5�O�8F+�(����{�bp��}��v����}�Ɵ����Q�9�� 굏A�zH����]���8L;zo{f�r��Oqkw-,/�R=��ٱ��`�|�zi�"3<j�4�#�k��wH���g�},��&!s�Wӕ@�qI<��ɤ�<��ҏE���Ք����R�%�?j���d���[�
-]HIimb%�C�T��/�U	�� �6&��i2��t�.�ۥ'�6LG�ڙ�"m�^�_�å3�|�J�\csTo� %��U�B J�bis'���~B\�b��I����w\�M�� r[D��tT�sP�xɋ;���.��VLI�E���m��H���;׭��f��9\�X��t���Ā�`�u;�s����B����,}����n	k�B]o%˹�4����I_[�	�6��"���o��Q��f7���������Wj�J� k�$-���9�T~���)Ӣ��0�x���6Ͽ�꽴J��]�'������*cH�C(7069U�f2���v�#�밚� �; �_T�p����[�r�G���p�D7{B�zE'�HZ��"�Ѹ*Yd�8�����v�`a�T(/��*��4)`~���%�zo�
����F�<݅�%*�ĭ������=��7��F ���Ɓc:���w4C�^ Y�eّz�VNjC�I:Պ�;"��H�����uK:fGޢE��Q鯴N ����e�;9a�5��g�-=6"�UGL�#�Z$�Q�)�6̗h�+�Q���&a�x�$ �	a������B�g�pV������i$'tB�(d3�J�k�Q�o߳\���`��q���Ɓ���&}��P��%>�r=������E���oʬHw���pJ�ǋ@Y:{ecf�GZnx��|��Y`v@[�,hM��X�J�9�[o�M��첫9]`�j�]�.��G��ѫz� ���^�%��� y�����7��fZix?I��Tu%+.���崠�ՔH;$�j����ŽF��?i}���?����A�\�&�̲N3���4�Ց��F
xȆ��'��������hN(�fsok��ެ=g?!�`�䳑��N��� ����)9�69�|HK� �?���5Q�Y�Q�����׵��'q����6�D�W�?��ix�x���T2���l�%��C�p��&�N�>cb|7��lK��9(\�Jwfb��1��w^��q�l�#�ٚ�8e=<C()��n�*g�8V���v����e���Ĕb�]�3�\ܞ�-���R*C�&���6�Yf��TZl�b�mp1B_dڊϣ�w��mI��2�x(����Xy�_S�`̨\�U��[m�[�Ϧ&Pc�k������ |~@[���
�y�+,l��s$��;	�w�|�G<T(��!�ǱP0G�o�xFNA��~����P�b`	��Q	�3��LY��x�WG�b�OĦQ-�13F��w������o��{���������h�P6B2,��m�S�nǽ�tVEo&C�rC���BMy�����k(W����G
��Y�iJ�t����5���hb,3�f���s���D(�˗�F��I_L��4��F��\[� 2�|l[LOL��s���>�y�U4O�'E�]f٧+p1,w(����s�4��)��f�GY*�M*�R޵ݩyQ�Կ0��֍�ntK���ڨ��h+���[W������=�=~8Pr���s�p��_p��B�P)��Բ6b?zak� #m W�\*��ѣ��
��D���9ޥ"��Ҷ~�g����[ٚ@��}����q�Õ�O)&(s�'�Qe�����ߨ3?��Ec"\���{�*�O��٤�~�(;Ǜ�(��)�t���	k���u^їaz��+ 4I^`1.��g�r?�Б;I5���_��<��X�#
��U�VS�/��<�l^��V!��<�$�u�Vc&<+/!=|fL���xr�(� 3��j3���C��F��mS,�1kx�܀sgVtǡ��%�*�C{�t�-��;���|d!M��`����>�D�@��ѵ��]��Xs���zY�-�u��q�g���n�2�R�>�^�U`�év�C���������KČ��p��f�o��"f?+�_���x���#0�~.Y�#�l��d�{e!���
��R/��ӥ��{��t���|��^*�\�rv���Ơm	�P�����u�O��4�{�!��,.��m+8�t���mqP9��.~tR��F(~Ù���d�Ɲ��7�b)K�� ���;�ā�좡A��;�$�)Ң����@Z9~(?�U��6?�	�5�i����R�ޗJt���3�KЂn&Z����^�AU���O��>�YcKX�N�;eVQ��ɍ.z:n�PeP�u-%v��t��U����JQ�_�i��/,L�"��֝o����o�a�+��|z��+��n�<�2�H]��0px�b�T�T6��}(P&�zJv}�\�3Rć�����'N�� A��zT�hN���S�}����r�{8@�%i!�em���υ�Wq�2x��X8�q��*2�\h�K�Za��d��H�qS9Ͳ[�Pn%�"���pT����-�,<�=�"MR��^�D`0(yF��_��)E�b �O�	� �7��O��ʾ��Rw�c	V��T�nf&���YC����)(��Bv��]n�Q�P�����_���#�S��	��0ْ�G�	j~��,t�:J����Dľ�D	N�)/��ꋨ^��_�e��3�]B<H�F9��Gf�	E�A���f�ɶ�x	{��Qu�˄�_����~,~#�_�����՛�&��Zwn���.Yc<�u2Hb���h���o���_p�֑-P�y�]�׮�֜����b��i��[!�(c�)}�a��Z.OG?��9�ݿ�l"���N�� W��<㛜�|��N������6�|d=������ z`�p�I*+���<*4�P28��O�k�+x��D9UQ$���&���KEV)��'r&�&����>=ҏ�l�w*z-S!��%Ch@����^�Ϻ�C� �O%]��,B䡜��a�qQ��7#��}"
f���}��(�-8-��iT�(��M����s�LA� ���l��w�'m
j��MV¬�8�&­�xq���iA����V��N@ς]�=|ݵ���a>�m��.WE���2�/�S@�����8�7\)K��84�O��_b�|���J�fi`I���)c�Ů_?c5�Q�	���@Ef(���"� �*��`�e���V{�Ƥ�VIu��?Xڄ��$��էnO����1H4]]�>ƇM/���!*(>�T��%�y�)�f�2vf��S]���4�Ѥ�Ά�i,��ò]���q�()V�ӭ�-�zI��w�OG�=S""Ч���Tï(c���y�hi��i�!nC��~��MH�Vh��ZY`&g!^��%�#.��ի��Ӥ�3�ͯ	�?(�d̤Γ
?ܼ�L�h�tbU�����;�7�|�y���G�
7`�� *�=��G<>�b�08D�7W���t1��l+�F|�G�V9��DF)0��틚�l����Ƃ�QqP�rܛ |�@���g5D{~7ް�.UZT���~��.8�`��pB�i�UhB(��ϳm��r@����<Qކ�r��C~{O�_���Uh�s���u)��J�.���m���|S�%vm&�!+��"�,�O��iS�7y�ن�������ט��ǰ���Zn��T(��Zk;I�HaT��ܖ�0Ջi��ţ��]�c��78�D�����%�aB�F X��ًU ���}���#�21�JiI?�6�K�f#��O�,X�mHFx�����˘(��u�&%(�Dˉ�6�5@Vϲ[�W5><LH��c�W������En�P��������_��k�?$�&�L��~�o!��˹~Q�-_�G(#�tCd��C �����E��b]���7;C�,^�9�h�%�t�S��������#�"�����E A�#AJ���f���� ���/�f��f�F�\��]uӫ�x���ΈGZ��^�C ���p����f�W���ߔV�WZ�TԑO/��p�e��9���J�ek�߷��9���(�e�97��PKfuI�P��`dY%N��IXz�����)�^��6f�*�%���I-[��G���_
�����˹�
�e�3��O�;\��<��nE�dc�4p���LBr/��<��-�㵊������{Cd��:g�//��q���"� �J!h#�9+�f�vՕUD��a
��狤�8�x���⩫n*�M��	��8�$��<)�T�V��ɌsKTK#�����Jτ	�^/�}-�X�o�KBD�?��!�C��X�]\����a4���h�Ul�^^�Eӕ�CK��!�QS����>x��P�j��~E
x['c���Nj�Pߋ)˰ej�䩩n����w��+�)/�ȼ	F:���LGɲ���g��6րn��$�V���;���5dݶ��V*���̦�Xy�(V�,���a�4�~��G�?p".�,����Ο��k��b[�Y�L1B�$��v"�/���T�J�3�I�/�/�	��B������Ou `��6�����J�t�]Rު}zZF�p# C�,���
�oB(4
IFQ��w�|�΢��Q��Π��Yx~�:��&�=���'�JkfRNԪ�u����#�n9�
��Iyׁ��;�i��#/�/�7B��k�їR>^\�!UB$P�}/���{������O�H9��`���
oF� "�Ƈ@�	�i��b��_����χ]�;u�t�z�'����:M�3R_n����2^��(���I�3�Q�{�����Rr�{���'!�Se�)�>7'���d��>W�;2���FYZ0� _���)������޵�3��NN��jW� o��&��%g(1A��,��ψ�C��R^��-��j׈���ō�tT7�
r���@l��ּ�������~�7I]���go8��y�L"*OLvB\A�'�V(��X��
�52������Bns�d_�s�aSVn���j�ϔ
[�l����֛D)<CIok&��9�����S��4&��4���|��K�P����.��f���Ϟ͌��:��:�/'�Q��{����UR;uf���1�[�0�쒟;������@|�A�/Z�W>Q�|Ph���.q>��]��c�����e�m)�͹˒����F\��� )��f�P�>��=P�NETp��MHĉ��L�P�M�YV5j�U���H&
"&m>���k�yJ��X�6�W�����;>#����&�^}��"�!�d���Ma}+G����,e�uRk;=6ӆE6�Dŵ���7:�C�>�/ _#~U�ѶH������U��ˆ�P�$���!Fa!���x���r=b��,����B=�7YT�p��a��{$�$���0Ն�g�6$QL^�l��,�I�k��ݴ��o 0# ��:�/e��*W4�ɳ:[���f�Sl�%�O9F��p���!<TE>�U�i�ЅIa�Φ��-�v}��F�h���B��T^�@'��-|�����se�$���
nO�I	�*�ɧ�|�1�,��H@X�v����Cm��uF|����?d�L��:��,	�8���r��3j�����6�N�=��g�;�D]�P�ޙ���wݾ%EX�F�r{�����k�d��e����t2�P��2��}�0�$e�x�4�o�D5��m֐�_Y��2OHX�F��M�0?��|�9H��~^�V���L��>	<T����y��:�S�%3S�A��t�O:��^��zEb�������F��w��qO)=�����A�G�*zhv��^�u�xy�eǓ&8���B\ UE��rc�TwfF��e�>���2��&>���2�ə�|�hz#�J�R�P� ��NH�U�.b�O���b��8��2I�����yJ,bgh�ٚ���wP�����y0�"��B���o�z,j$rJx0�}�i5����
,cY�ON���(4��aP�(��[��M
h��j�P9�6!z\Wnu�2S�1ju�c��t1�X�G�9�5ǦH�\9B�ƂH���p�8{��PD��2IuL@?�c�Vġc]
z�nNS��vHE����֎�k#l��D�j)t�h��̭)���Cr*qZ�x�x\�3֮2-A9>���G�AX�&.t��;�K��7�A+7+コet���{����ݘ�б���@�զ��¸+j���KÆ�5"g��w".E�����h2�f��'�~�襻�N�ƻ�V��>�9D>b��y�t5�Q�9c�w�*p*�1E0|�����vǡ��V	������2�Y��{?4�^� Z:�(��?�2�����Ώ��ǋ�;5J�e�><�Q� fr�b6����$�d�wx��׶^E���A�=C����"r����H熾�9�B�����+V�&�����rBﱐ��`\c`8F^��<A�X�2UJ='R�yj+J��z���%���i�E`�tA@^-z���`��;� b�	�0Ul6�%���W�yg~C�>zY&�]:Cc_ۿ2�^#`ᶒ~�I=*T}�FB$�{Z��v�nsj�O���q�e 	+�ީ{�i�p�"��Nǵ�k�w�JmPK�@xB�H����.R��'�i=���i�U��k�왌s����Y��yC��x[+�1�k �]n3�wi��Ah�',�f'f�+�$��WT7p(�)\��YV�]i.	�F�K�9_>�.�ROFB��p��4aAc�S�%0��t�5&�ʖ��w|�����_���x���� S�ܝ=\:b�Jq�V�Am>�(�&����ed^3G{���i��y�R��vm�O�*I���J9��e�+�o+{>.(�m'�b����k�S46�^�5����nx#�詛����h���t))|Ě����q�Z^ `+%u��t�|�d����"F�T��L�� %���~�T7& 29X�����ޑ61*��}��)��
/�9�������4m=��o��Z�V�d��غ
�ǋ"��?CU�h.awl�v
){�rǇۑ	�tJ���*�L-��`5:�R��|�#~L�:j��t��)�N�kd<����i�����-|>�*�qM�!���| \Ms��$\||�m�wX!;D���9�Y��T���&Y˙�O�A�V�Y�����k���U_���0+�]�g���q/{8ToP���	�-��5��s�����j�rB/�����H
��^���m$d�8v�������g߭�տ@��ػ�$'����	�)M���;�7/��y�H�ȕiK$(�=%0�������s���I��l�kK��1�Ū�D��=\�I.�zLw~g������|i�xs����)��ӓ�!�D]3��e��]�!O[�kX1
.��P�T����Ԃ0 '���t!���wH� g|�H��<��[�
q$��r��/�D�1X��-��������-=�v��eӎ�\��#Q���d�1�;��C���f�M��9�)I���#᳷��R�[q~�%Ǜ!����~��n�K/��T��#Nz��nAKd�0r ���P�5� ?��W����� `��Q��0������� ������D6�::�j�pHAt�u�qg�bb�F�[�9ST �{�0�V���H-���[� �.������N�"����� �ߍ���{��N�5��]Xr_ZKs�ǁ�H�V��N� ����V��da�9��j�Rɯ���"�L��g<,G{��c�*��Q\
�nEHվ�Pg�k�n^���!��	#(��6�ԚR]cS�������f�z���7�
�o�4���!�Ny�B�>�:�~Ѵ�B���v�12nM]��m��e[yE��|��R2���gZ�-�..�Z�����n������L��ź�o�޽��51J����Xv����Z�d�z|M;� �&&��p)�/Zt�hٺ,�d$��E�\�Ra*�`2���՘�K��U����#m�ٜ;�9���
)��8/����Zp4G`�)�с,��"�Q�\�Zb�y�x {����k��dAR����j�V��r���UxL]�MĆ�գ�^�H�p(�b�ޠ��LX"c���{7.�����;�����"/��E�}E�q��(�ʛ]n��۽���({|ʤ6�K�0�C�CL����d���tW\u��Lub_���(9	DF}C�*c.�	�W���|P��/K�`k�@����#u�:�����+aeS�J��fXH��D��?m�W�ɵ��KL৸�I��ȕ,�/�(������O��>�� ��i]����B��ٽ3��=�̀v�1���zt���\�0a������!b��k�1�N}���{��]_lPQ�6�V�NӖ���:���F��w�L}K���c��#�����Fw9��<� � �%0��#Z�����Y��_��=ا�F�P������
K}!;O�����U�twz�r��/��a��[���v�@q%oYG	���^``��"OX�@)S.�t��g3�0�ip[��/n�;]`��	�S�?S߂N{���_�g�I��S�܁Bz+ݭ������d�y�aKq�N��WP���&r���D�~�������{���"0A�2���3ͪ���X\�_��$�١8���EݙS�y�$l�<�V�_�y=�i^�9�gY�&�~�<��ǣO0Ú����4�V�LϘ�%�e�z���W�W�@P�������Ɣ\��[>/ݹ�"p�e��c9l�{� �<Z<s$�t�LȻ�30��J/~����M�/"sO�r�&X?���{����]�������y�P����K�`[c��,��X}�t%s#k]O�psjM���Ya^&��F�lŎg��2��َ��݌���H���o��Q�2�{\k'?�e'��0�/Q\Y�Js��3p�?oׁ�ME	��PX���ɭ����gLᄋ�7�0Ρ4���\�b�#g���}���m$�/��Z����ך�$I�r�@%Q��pJ��	����t�aΙ�2q���$��ha�r�g7��6�+
G�U1t��S$�����Q�$e���ǉ3*�:?R&3-?�byXQ$x���4w�޿B l�����^9����W�u5��;���B�=☬�ݺ�~u�ե��T9�1�4�9I�GQ	�d7�����&��;D�>�Px�`O��	ϴ����w��1�*�&U���ʘ5�`�
e{��.6��0�wK x*��$"��N�Nzߏ��a���rN�6�h�� ^�|p�����Ǹd��kkm�=����kM��Xl�n�\pE����,�#�Jz.������:�@������@}�s���}�B���@)5گ��¡���y�e��y���"�RR�;�L2Xp��sG���ZS���ˢ��s�n�Q���Y��|%$��H}�"G���ɋFP/}l^!����c]|��8�;"Ȟt���/i[{��%�/&=p��[[���1|A
��j`�t���0�(�wY��,�%8��;��b�l�2p&�|٭A�m�w)�\�z��S��9�TB+g@�X#�~�Hv*���T%i/VQĸ���<#d,@G�Ӝ���Ȋ���뒣�?֏ڏ���ZA���@���i��7���UWǱP�b(�P�XiK��.�~�廛ߘb٤�aF�QU�r�ݻ�{���$�]�{���TԤ/���7�ӟϾ`A0�N���Ĳ�D��`���N�o�V��W[J➙ba����)ݿ�O�%�z�"E�0@�r��I=n��;g.k��+-�ɛ��$a#�z��#����V%����D�c� �Iv�r�'�_b���"��}��F�[)NK"��ѹ'��F2�M��M�Y�Kbu�g��[K��R
0�E����q��C��P��և���z�H	t[�<��not�࡜��	Kx�BEfM���I����� K<���ث�8����4ӭ_TFxs��uQ�ʉ�@�1�>����).Ǖ�ZC:T�L��u��XM�R0���Y;�9�\5&?�Ulו���
�h�7S
G��vU�?ktm?\�m`*f�N��@t�ܥI�{�Ū�X�ylb�n������<��$}+1am�cw��8�9�27�N�� ;_������U��i'1�?�(vɯk|�|�`'�m�՚!^R�O�$��X��G��ؿ�� %�(@�9�� w�D5ɠU"V�3�;0�R�E���0�݁�Zp�ȚXM�m��j.r
�+�ZXi 9>xLΉN_�ߣ &���u3�v�oM���"#�9rꌨs��@o���f@D�k�����VY�N���P�����	��Ͻ�p����&`%�t���c�ѫ�e���%������/n��X��`¯���`F�ύQCj��s� �I|m>�4Ⲿ6��n�9R{�v�lЅ�:p3ip7�!�&
;4��y:���"A�w���*�LP2���5a�CmaJ�\[�o�Z�{����Υ#s�1�8 ~�L2��w�3~�E[����A����{u��v��B�j`��e���b�L���O�/}z`)�-��B���"R��snFT�a�:���i^b"`?$v�㝩��]�zW�� V��w�eC5[Ǎ�]��b��!�V%��g^��DAN�|i��c��R%U�Cx���O��sw���1/�m�k��N�<��|�0��qz�D��k/������3�eOg��G��r��B!��ϸ���y�r�t���y6���PQ|0���;���Y勤\�� ��7A�3h�����Q=.���R~c8~�%�������x�2Y�X�-z;��2e�dh,K�:;�$�ȼ�g`�QfP^K99�{��	��ɟ�����!��JIL��j��·�D���֨?��CvЩIz�3���O~���P���3�.z����X� N��@#��L�l}����:�r��"뱏�������X񓫞1�|G��@P��2�Fk�O������g6��n��k�=�i���(�u�t��&��O��v=t�Ĩ�Cy�2m�!wr��J��[�+�w��~3j��V��'Q]v�s=JO�	6����v�:pl�0G:3���tK��[�DpY���Pc�<��١��N�k�>��n����56�$j�(�S�)5����ev�W`�g���k�q'��e(��h�>w����0 �6�Vn`��w�½f"��2��TV�غ06ٍ�!/�n����R�Ƴ��A4"�ׇK g��}���j�ʮ�K	���4J�ѷ�������Jf}�#=��(���j�1=f4�8ȝ���Z�L��K=V�.mPۇ^�7�jZc\�G���:9����v&SQj�ah;�+�#����U��Zi1�I2?;��� ����`�ȕ%FP�����Yĉ��m�!uÇn�s��������_�e��"q��v�����N��8:`��\G��Fa����G�	J\��
.���U��`=�F�Jҕ����+`���
b%,]��a�e8ݿ�t���f�-�v�p�]pxߦ�r���EΙ�������GlU`mHA��[6����R�dj���&�j)c}䭅�=��k������7� ?
��5�Bi��~�1Z"L�g,��3���|{K:l�?�th�e$���$�	$����y���E,�����_��Z��UC8	j�?�ZQd�F-ƾ1�O��E�̞DU^[���Ɣd�\n��	�Ҋ<<�s����00�+��C��ҏvB";��(��  }�h����Kѫ��>X�i���+?��l����.�&h�g=�:KX(Z�S�a����y�@��$�r� ��?E�׃�<��|�����<���k�IZ�yk	��<�zQm�a���?!w�s��t��o�Z�>��z�-,;�A}9�C�ɠMh����1��g,
�.3w� CY�/\�*�b�FB�2�LI>���f��Gq�;@n|���g�f�E ��	�a���8a���`xfC�$h�O��"g�0j���íy��m�?��wT֭a��71�vJ�,:�X7sdd�k�B4�p/B�LF�����3_�T�[�D3�ώ0e�����*�Ծ E'�#׭Ew:��@D	9��^�9�q1W׳��?L&�HW�x�T��ʊ ςl�V���.g�!u j�4���@�o�D�]k��+����0��fhՁg=fq�:�sI��U��n��1��	_
����r\����w�lDҷ�Tޢ�V�54S������!�I�mc˰����u(��M�x���7\1�X?�Ύ�?e\3�9r�$X��:=�0H�`D���(q����v�$��Z ��+خ��B��[Q��㵿�њG���,Kһ�,Ɔ06��y�U�ҡ�8[IGmj�\���&�*&�:vYe�$H�ƌ�����&݊3���s"��I��c��H�WoD����RJ�h�S��z�hO����D�W�c�I��`	d�s�z)�N(Ѐ�	Д�{�/�J�F+��Dв^Z|SzOvb�E<n���6�̟���ƚ��Gg��z�:s$���1W��M�9ږ�0�ЧM>�� K�b��R���%��B)��;#o��Y��xV�_s�k�dޏ��o�У�g�A�����К�1���r03ݬ��7�mD	^�5���/�YLUgw��.G�Zs"vrVM�'�K�^X��>t���~4��y�ư7*5�$<B��qv-4�/�[5%���HT2����߷���QRSH��N�\�Y�k^�E��o0�l*���`�*n�m�#QZe���I\I1��<�M�J���6�sA$\;�)Ћ��ß��u]�H	����˥� �4�`������fH\#�?�c|	4������Yh���"ہn�ۦj�s-!KB%��D�T�8V�����뼼˹5ws�Ň��������9��n@�q�Sⰱ�m2"�Y߱�e��ԫ�	���\�o��]�Ű�w��3�X2�j�JK+-� g&�90��������[�[@t�����})��l�e���܂Q����J��H-Zf�AD�2��[ww1��Z�o��fٳ� m	7-���ψ��9+]k^���AJ�q�OPK��S������8�^˼��e
�聪�Ys:rq��d���gƎ�]-S������z�a��#Y����4Y������4����2,PG_g�ˑ޹q������[��~;T�Z>��J�!z�J�?A⌀XǓY_�`j�{�����^�����j��L�DpsK���3ˆ�*�u��2@�;̋�C"7��k���;������y��X3�/j���zM.p:��]���pr�!/(ה֫1WZ�zV��A�D�T���'[C�۩	�(�PX��S������?�����<J=歹���Z�Gi,v�g�ͯu8o�r�����*��[�����A�dmas�>��2�@vw*�iP�}#`��J-A�KP �I�ڂ�%�扻A��@�N��hŧ$x��k�:Vi@t���+qn��G�؅
5/�����u2�8�!��a��'�h�!����[��k��ݝ��y���!
�>X%�.q�I�T�8-�6�u��)=�f���<�������b{�F��J�"<D�����A�*�6��ia�P���|nON&��)܇4X�x�Ҏ-��)���5�Zhd���`R��q�����@�嘗I~�%�������yR��B^u�%,Hz�!m��lM��ח-$q����q��P������o���η)_s;�oh��W�n�u�4[��������C�1��	K�!��o�q��(HZ
��v�89�T^����N@��ѡ��>�a��:�C�k�K?�Q�d|j�����%��)̖�H��i���a��ri�!���4N��X�%8�e����8�D��È<*��������N!��n�A�6��h}hwJ1-� ����I��Z�~�����]���hD}��j�"?�ÈѾ�{�C��Ю�l2�H�����N݌�mc=9����o�ӥ�C�y?@���g��~��G��͟n
N!��L��eUyiJ��0'�řc-���n�QC��������J鑡
��":l�&�k�ˠ_/C&=��1Xh{�F�~>���g'����9Z:��9.>�B�-e��Eu�M������瓓����UAGAUȳ�3
,�A;b(�s�/�gj���rv C�ѵLj��F�3X'vS0e8K��r�H]�ٽMvК)�H�?U"a�48m���@�����>�U�����-Y�I.- �[r��+j�݋sB!8��Fn���H�8�e���ag�<����lS�.;�C�'��3�40�֦в8�ѷ�ࡘ��;%t��|57hT�kY�N��*n�fMs3�`��y���/��ՈxE^�����W�}�� ������m���P����o6;�=������,-�v�`8�D KQ�&�@8��`��툃���8�{��
A���`C���)��0'eMOI�u7��
.�"���Rq�"�F2�)}����v����i�o%م2��>���Õ�ї�F2���\P}�J/������h���ʌPQ\���&OG^������[H �ǜ�nvȲ9zY��	�N�K��F(Z�u�ׅ%��q����?���S�{3�/8�=L��˂�Î�?LS�9�F*O��ϳ�?ȃR0[<O�R 1[[p����GmŸ��3]j�e@��W� �v.�܄&��K�5��<O�}���a�h�������_6�#:5��LNH��qfy,�BhV��&�T,j���b�#cdVse���-���j��e�J�[�f�H��]�D��{�Õ��P#^{cg̳K�m�P��/��cwJ��h���w��p�M"w�>�G��'8FVU2 @��l鏢,�י���D�� �p�a)���C�hD� �	|	OTyBhzq�8��N(H��m��wK eI�<f^B�&�t�`�ϵB!��D>�lj�->����(�F�\*
���I�:Z�v��?U">��%bH��/)�z[|�H¦�J8�g�?�uyf��	9c���'y'�ث���Qs��/\-23?�"/�=�+��l+8Y��C�<����*h���D�̦N�A����li�urT��"&��A���.dO9o���U�a�r���9��-�)S��DO�֚���Rā6�x��,s5�K\���WVݮ���C�K^�/e#�u	��|��^���G-A3��ke>NG(y��^`G5|��I]0�v�����ުH��vh� k�h�꿋��ڦ�4�3m��Y�tnw)���7��}R����Y6��m�Г}�$$�ݯu�=��R�{���s#���i�&pf����܍����	����A��(����f3��ɳ���'>�n��e�Eɗ�(M�� +<����	���DOˎ��"�,�?nŀ��'Y_\�Z�����#���b~�������V� lb{�P����ެ�<Ͽ��� 7��N؇��3-�A��@TS��ePL�����1�V:�pĩ������;�b&�|�,�u���W��I|}�
W�u���aߝN��:�SpYz��;�_��U[~�s�	�G\���Q;��i�d��E�i�?i��-� v�2�W�����`by�~�hC�X���8uB�v�͕/��G_nqv�EB��<\dy�E�pWV�gR�ͿZ�?�G=���͠,����?a!�~WU�9���<R0'�S����p�'��a �pƉ	7GM�����i��u�:r
�ldη��s�V�n}jῒ���.�a�k����Aq�ҧ��Z�Wu�)(� >-����vga�� u΅��Ϯ!ʧ��Q N�V&|d�ȿ�x{���B�.B�)���ÓRBp��ZY��7���00A�m������N���]�{%A�SE�Ŏ,���X��^��P�gYu̓ ;/��j���]#�(2[�;JEǣ`��w�b�W�E�$id=�A��&jn�3����N�!��fL�/ɳ����,�o�ǟU����?ocV��k����y���E��y��Zi;���Y�d� FX'؏O�#��2�.�Į�-nFe�y�*�q��e4�w��0��q��Ǒ��*��^~�-X�M�F��^,������d�M�/y����]��V��õ���F��da� �(�XJ��_� Vd�+3vȎ��4���M�,������uV=/�M5�"�[΂��'�z�6�-����D�G��Ώ�p�i�}4,�9�kl�H��Ձ�f�D�.��-X��_��qt�B�#��GW�잭T]6���<(���+Xl���3�
�$^jx��'YY�u�"�D-쓟s ��S�4����n/�)�S&��0�aw�r�H�J�e$9����KJ�i8)�O_{U��v�Of��0�.�M���% ��̙��鶤���`8_tw 1�I�I>e�з��W �ͣj��m� �F����V�V<�8e��{r�c��wN?�6`2��]X'���p���;�O�m��P},�����g_RZJ��,��a������U2�҄o$���F�ߒ(��ү9��Ԣ��E�Q$�6.��\�G���������bbs�w0��5>�e��$��\�+�
� ��M5)]%}�D9�@�Βۮ�1͓���zhnO�݄92n�����r��b��?Vh�����8�̮�p���0�����a<p)�'��t���d,��&�ݾa(�ꋎ�G�*[����:;8;�hK#�W+���!���^e�3���դW�M���2ᱭ�i��z��7�k[J�aL͏QZߚ��W��K�Rg��w�h�}q�f����]W���/"$k�B@��(6�Kk�j�9��B�a�˖�f=�\J�Ń�4�۶�HT�1	�I7�}�Ek��lf�Q��/;Ȣ�K3=2lu	6[P6e�{Ԓ�)�3$�p쉴�!�J���*Fu��eg�۟$PoV����Ob���b`��:���!�\�����z�Q:�^
��~�o�Z�ә���=���߬�e���	�bI�(�:�Ӷ�X�����XN`�8C��`o9��w�>�wl�yP
�{��~�D!B�-���"w�{"�}"W\�͸7^���;d���i�r�xQ}���"�
�����~��e��B܀,��I7p���| ��-�S��!�{�	�EW���7:��B�P�
��=&V��>��?����"�}�au�TJ��f�](�e���ULU9"X�L��Ѣ�/��8��Yw^��S2�%lL�.r���_S��ˣ�A�P���>�8z�	6.X
��dϸZ	NaCZ:�Eh�!�?�Mb�5�D����#�ؑB�n�؜�0q�����'�1�X�HcS�e�Y�Hg���VA��l�_�n%�l�9����H` ���(��BL�O�Ӂ�R� �/��d����o�*�����{:����B�m�'���{c�`I8�_���;�|:q2��	E�HK���)�"�K���O�+te����;�5қ#}L��j��f-�@[���˕e�J�1�-��r0|�`�5B�p�d�xQ�6��zF��-4���V�z93@킂����=���6��� �B ��1��P�;������Qv�T��&G�%%�jc'S�n��^�^�w���[����lVPH�0�{K8j���	d�.]�Ō:C���h�J{�y(as��_��?`�8	�~nc�4�_���;��1S���Y7��.���� �����o�R��n�W>���Gs����TdH�+lt�i�J��K
ow;H3h���:xG�M2�\Y����s�KpTf]������"��F��S�A���O�`j�yp�.�5���1��r�ٿ�z~�n��>�/�TvH�A9%Y���1ɦ���On�陭�j,o��i?!z�$�4pG|�0j�t�gݩ�I�����!����=O�XL�HDә�S?ǭ+u4�31��T��|���On�\�ʺz��"��UQx0+k@��|Ng�6������ZMB�\��u$e�w���`]Lu7ٞ���������z���/� ��)�+�0&$6؊@���A�4��b����F[�����ϯF���T^�2èטy���ޛ�		��������jO����R۫F�0_b������t.���,Zv#�j����h/���I�?�9����՚\w��$L�<�3�@}J�ނ<�wu�(��r�<0Fgk��ω�Y�W�~dm�%	\ �[uR:f!������B,�d�9��F=���:���Tv	�zLBC���C�dh��b��V~ę�ӥ���!�^F`H`�-J���B炁"�η��|��?�׾�Q+�z�(�ὑ�`,F/jH�mi�Z|�[ZC΂^�ל����fc�P��J�*��I��j�5��W�y|J����ș����<5îی��ў˥c�ܝ�"O���*U%��y�?`@����D����έ.6s;��_�f.K&������=ν%�bPg_!p �'���FzWg����ҁ)L�58ܩ���T(N7��7��	4��)R���@��[�D���wm)Z���$� 4`�9r���r-�7�	Ch2���{�8h<��V���v"\2�5��=� ׏�A�(v�B����|�]��e�+"i�7�Y,g�Rޮ���<D��*k��d�䁘��d7�Zf��U�-RΙ��n������}rԏ8@���BK ���n%!0�/Q�-d!���:�.����TYV���ʉ�!�᪀făiJD��2�m���8��)���F9ۍK�$��0S6Sl:T��h�����E��7d��M\�����<~�t����^5�\�l�4��P�!��� ���=�����ӯᔝצa�W؅�Lc�~"L����� �{q[:�u����$�ڮ����t4{C���鿿x��D]@[�;Ǵ��?��K��=C�:ܤEWє�ģ�>ZZpn6ق>����$ȥ����m����v~��^�D�x }7'����T���Bպ��)��X#����ݛ�v�9�p�ǆ/L!:G_��|�r/���K@{e�Y��@��&�&�9r}��+�/I�{n�a�\�͕ɮv��T^��k����9�]���~��\Ug	�!8��q?� �������=�yL�������f:�?��!ބ���rL��ҡ��*�Ob�rs �ٗ#
a%��W�A���2�ۊ����o� �
������LZX,R]*z�^489k�4���D�%]�C��EI,X��߅"�c>�"J�r����%��בD�u��S���,b�NFM������Fˤۉ߯�z7~��$�⸟�����z9U
㤜h5~����o��"H��.6{�-)��(=�]��D�c$L�u
�_��VCj܎��K�Gzj
��?%��~su���}�""'TFK��傂���RK���v�ƚ����r�A�C��{��v鍱���\٢P�g%�%kو��{�D>
݋�@�����C��g��Sm�Rj=	{k�s��@"B�M߆�=���=���*]�9�䢛>����悾��� ч�������c���B�d�(	���Ll�T��4��a�R1�N�u�q�p�k|�����FRS]�;��� �
�ྐ��6l�Ò--�����Z�Ag.�S����.��;��Aѓ4��h��4��*��D<f�()f������}��rXE���f����½S��Z���J��}s�L����J	���xR4e+ͤ����g�dA��yWp�<������\|�x�I	$
G
[8��J���tXK����'�ZA�D�+�]n��ȵ<���,�l����ݛ�~w1���Y��!�Gm��Ɲ�F>��q{���'iZ�f[��5_���΢�D"81��S����32S�d�0	i�7��؟\���s�A�ɖ�"��ٜV�.ܹ��<��/إ}n��W,��~wfݵ�p���UƬO�p���u�R�e�AS-`t����pB(��L�CCp�����2C���������:JD��UWw��{�s������)Ʌ3��S�0.����;�k�+��G�0]�������!�ԑVP��u����: W�����'m�W��T�h���my<� �R'`A��R�$&��L!�/��b^��.e=/�z)ڐ�+!��~9V��V�E8zo@�6�;����J��e�����T������=xrW����_ǝO�*� �RdJ`��5����:�y�1T�����֑r)n�k�ݜ Dq�U"n�!A�����~4gBq�u7z��������E(�{���ڡ+a7"�+���Ή���?Z_�㵤��X��T"z�����{���� :�<��=Il�lOXt�h�B��������y^�I�����!U��t��V鋰3��#X���MgP��(�ذd|;<��Q�>N���b��q7G%��+~��uA>	��n�R��&:O�#AcP�����Ap��Fo�'dO^A�~7z�|\���ܖ����H�-�+۬VQ��)6 �������� �U@�&�X:B��]~��Hq�:�P�fz��R���5�E� D�	�|����s�d���k�������{i�DKz��Ķ�AU�X��^���^dT�?_O`�"ϙ�޼��E;�y�;�qL�
R"iwa�â�h$jkyZ<&�'z|U$�2��S�
��q:E�� �����?��-� ��o:��j���~U�/�&8�g��"��L��a ��o��aS�+Spop�&�<�8>�ЬB�i�:v�##4��w��<��S	@����H,yDM6S�'���y�őm����Q�?�&"��k�яX�g�h
<n�֚هwF��w�^�ǿ�^��%�z�u�)�	�,q�:���)vHcK�GK������1�|&��N!�6���iʑ��h�<|9��+D��Κ�֐Ļ���)Mx�>}�]1@�Pf�����QN&�Y29� ����*c��mQ�c�J_�/OM�����N*����nuŤ��/⑋k	��y���v�d2�R��f� �yp��I���O�(���t������ް��6��Z���'��*����*��Օ�'���
<�{�
��+�?6Ea��c�k1��fL1�����
���Ƞ�ʄd��E��/�&%(����w]���2&z�1Xb.A��hu'm�!έ�Jj-�j���$����1����9K���[�#^&Hė�ؒ�c/�6�Y���l��6%�q~�Ѽ�Е�3�h"Tft�I?Ҍ"Pt��X��C �����������[ʼA�㇬oK!�I�NW�n:��E��)��w�W]��0\�H�Ŷ����¼��b��x��F�\���l�L�N�m@'X��ҏ�GF��KO�PƬA�����x b���쁊��E'�C���;D���~ѷ�(a�����˿��k�YG���-���$�n9��=��d�;�b�tB;tC�66ԄYW�7ʦĦ��_�3��M?���7�����9>Lk{�+v�����(#wƠ���VC|���B�$�,�#^F6�s��E=UsR��Qpom�Y4�;�Ӌ�07jcC@O��}Li|u[��XTZ���םխ����|� �#X5��z&1���#������&!���o��Ý�,�y:��� ⡵�5^��z�}�^���t��JeZ�Ntk��%����ҢY;�3�B.f��y�.m}���n�cl�WƒȲs�h< �����$�"BhY��p��@P��pŏu�w��;�g�>����졜��M��-�ǋ��j�חNM����=P���]mXȱ��+ls�Q�f��<Ǿ?���M7������u;T���3v�Ӂ/2�j
T�&���;�g��7�]�N��G���F��-�/�����?x� Dh��Y�%L�랋�
�g䦆2�pEI|\��.�r��¯��R7�53&�&m�������1� 
������7e�f��W�?X�o��e�J���U�'7�33*�1|�]���Ei�^��]��P�(ݬQ)<$>��� ���b��aAk��s�T���j>Q�]��5vV�� �����?IܷFTk�8
�sp72�lO�%_� ���JT�'���N����
0u箷�mA�r6�}�籖���o�ҋQ��$(	0�����Z1h'O�9[kBiA*�s�]�D��c�?��[J�S� �������ue�EIC�c�A�q�j��(k�(�+n�K�Ō_ ��Y���5�0X�d����5ч�&�����M�u_�~`cF�[�4��J֒�`�xwt\�/_�U�0g�;� h[�(����U�N^5�&������6���L��N�|�����C��-kLI���J��e��%��~'@Q���Z�hU1�, n��A��c��!T��E�����'y��*Ѯ_���}U�8�ہp~�Q�PƋb��^	��!ZmV�����vY/���9m5�:���\�b��7[�/��?�[���À=��/�� A\P*0����i��S��
���\l
zw�x�e��Jo�3c��tMr��d*��;g�_X�ΚV��&&�P�h��Ip��̐�������v�3���E�~���˹��l���5#����Y�)#X���A"m�b{3(��������E��t=q��1�h�A5=�� u8�P��T\�%�T�-x?M9_�D�Þ��"Z8���x�=��� F �U����4�t��ۄW/~Ĵ������bXƮ���R"lD�'���h�)T�I����&��W��§�>�o*�����Ke"�������\�n�N�E�o�&��L�]9�NL��K$�_������Ĩ	���1����VOp&-^P��Owpe���|BC�%o_\<��?	���G�+Ha�m�2��s����k��>vE�!�kȕ|�2�r�����6�r�\ �˺_zm�5���F��x������dwB��`nή��zl��%؜�;��xɏ�T����\����0b#��4�!<R�V]s�*r�O%B'�C0A���.��܋�?3�j`Ɠu�%ge����~��t��R饬#������e���������|�Y�_�S!�5��8�!o/���-0��~7Q�A@Ϲ�I�C��O%�,q��?��טW�0׌ȥ��J�k5�g7���:���{��ZU�������˄� Ġ+����S�s��&���	8؏1�w�JҒ�V}A��&�<���#��i���fe"�?�����Z0\�N<�>�~~Y��v�S�2�=�v.��66�@��o,yL!"35��s���G�=u���k(�	 �'NH���َ�D�D�;����I�5��5�,��{���Nz���h ���-7�,r��$�&N:�gwvi�.�蛫�B��:m 
Y�?��'���x�ʊ� 񃇉r�� Y@�0~������jd�.��3�ry?�&�ؚPyZ��hN�k}5C�^+�̫�����f�Ni�)����b�>�ვ|���.E+�; ̇�	#D+��O�ޗ�UC�i#nȻ����3S�Hz͸����H� �:���O��Q�H�I`��λ�~χ���]�Ĳ 6KR�)���^�xX���jF��v���7�������BY>�&��1� ^ER��D�^u�f١�&�rv���P-�r��x��o�|0ޞQ9<�� LotԪ��hB]�_Bf����E��T� �G���o�JG)�h�>gXSps�ݷ��롆��Nn�� )�P��6��~=��X�"���3H�&�=0����&\olSp�ܿ�v����	���0e#��$��J::^,捘d٘եҶFư<�,�=rV�u��6.꼭ɟ�Q��{,J�0 MF~q��S����錙ڋ���*�NU���w�N����Q�����bq�^��6��'TژR�mĖ�rf���X$]Z��&�6[��������L�Mg�@�}!�d�r�:�l� ��{5��]xK��WS"�jcŮA�q�\� �'F(��V���l�^+θ��a�����r��hNY@]o��������"�8U$�`�@��9�L�Ŋ��юp
���5���e2f��S2�I�N��&�n��aY��J�x�}έq�E�Z�]���hﺦ�v{���K�M�� �?z��?@�a4	�
$�^���B��?� ���U��"�����˸NJ�����#Qf��.�	��k��O��f��R��l��Ün�>\ӑ��}���+|�{�k`d���*^O�ߒ?� ��U�����{o��J���ѭ�JBa���p��|C?�jkж%Xh��m��8�K+��90ڸ~=b��Ӭ�	"I����M��MtƗi�{�>LI@����,O��(���%�xO���?'����V&M��p&��FkAh�/Pq�����˚��j���j��r����<0�D���|j�v�^x�CĖ���-#U�e�Ky��v��8�k���ؾsy:���g:6�{��'�đ@bp f�^�'N{�5Y�*�#�ma�-LVC��|�}�����WU�f�Z�(�4�4�9!�����)��'�~�<(N�V�W�\���b'F0υ����kC�/�-�}���/�����j��Kd�eVb7�-��Fޓ���7*<X�3�Ьϐ1�Ag��tXFՉ2)�^&K��Z���J��̈́�o��	^0���Po~i��cF�4n�kB�L�����j��5s�^wKI"½�M��C�xS-���wq������}�U��`�z��4[�����z,�9�`UR�2����"�1��Ôop~1�Nu;d�+��y~M4�`N=��DA�B�����N��U�DZ�b�Q�u���S���|u��kwq-VK%�s�R@۟JP���e�t���A�����?N��M2a(��V7}0�9}�1�F������N[������8r"GC�DF���@-��|�ͦj�#n��g<���C���=��j�]���,��  g��*��I����A���p�UM`��E��D(�,�@�t���~��������>�	I���Ll��n?�ܹ��?�}�ŉ�����m:����L��/E�Q#���9�a�:����Յ���8ƍG��:��a6wz���=x�{����>�y��� � _i.��$q��|�<v�=y��� ��Lay��-c��`�׸�J�sCZ<<���zB_�`���7$��k��DJ}}�`��>�GO_Mخ#���J�u�x��7�i� (rD&�U�����Yf�dy�� 0~�	������"cȅ��W�]����I<���t�G���I�C�s((%��N7�?/c��̉i���^��+u�������O�-Ȱ�9�o&�ގ�/�+�{�~fၪ��v擉L�t��������ꪨ�P'_B��n�_��<�&�������u���a�1�0=(b�|�r�s����Yi7�}����ߜhw����i�����9�!Gڏ�N��A^z�O�<�{�'�%3{8�i'ۗ��܏��$lYW,?�U5W�q�F�[��˱��:Yz=A�~ͷ �5�埂;�̍����+�h����qʜ�Y�UI��Y�|A�ͣbk�j��tGV�^�_���h�_nrzƣ���:��+-��%��j�����V,�k-�҇�i�[�Q�đ������>�Lyʺ9��v�9��a�.��%رtgZ}�Q�R
Oh􌍫����|w�<�aۅ�
H��	@E��)@u.�s]j���5��5c��2s1�`��	<^� �%r����o�g�6��0��̢%��ة8���3\��Y���OcX��ed�ᘜ!-��l�J��mJ=P�݊���C���cq�'Hp�ӻBPE3�x��4ϕ�SP��}��Ӕ7��m@��J&_l3s z���i��=��~#JVW?�o�̰��B���1�T�}ܫ	!���u)	՜,�y"��������!(.�mC�l4>�EX� �j�о J�N-̛i�����H�~)w[���m4Eϑ��'.�����洡x]��p!��2���Xv�b�әVJ�|�\Zm,�$x�x��yZ4��C��e�6�Ƥ����\ɚ����֩8��`gp`�u�~>�ml0�B:ߙ�<�-�B����9�z��wn7� +����ү��5�|P&YH�,���_��սuRD'd��|�0�8��&\��Ѧ���KM�P���)K�� �<)=9y%�����"�������I69\2��	���xh����o�{T\��dz����B0Ѿ���Fݯb6�f�����1q�����|�po���fLv�Č���;������vLN]��?��FZ���B���(�����
T�_�paŶ��>��*m������E_Sk?�S�m*g�|ׂ�}�Ǡm6#�]B��l"��'�����,�=e?��>L$���Lo�"�B���2�2����r�����n�ma��r�)"9��UD*�	��ݻT5q�l��g*�K1"�fF�ĚF���O`1m��7��89�^b���B���:�?o@DCk�	n��:G/O�Ɏ���29;�GnMX]��J�?�xX�))�bV�V���n``J�a/\A�C�j�A`���V�=����@ˁc�O�mְK�H�A&����$i��h���"s,i7{����wBQz�BΓ��@9.x\R/�c:��B��� �?��@q�O�����ϴa?��^��%b9��I�}ZA�@��ˇQ�4���9�gJ]�}��%l����ʄ�|��u��CںH��'UnGRY��7����L���R�v�bEw>f����6���J�ҹ�
p� qK?+����"f����Ӆ�����-[���x�&���;�t.>Y�e���z�W�N+��E�(�=Q�U[���/
w�������L�����K��[��)5�X��J(ԋ>�#l�8�Dv�kE(!"��C	�B������m�ۅPL�<m j�z�-�HSc����W�t�H�v�&��V�	������p*Ғ��e�ڀ�k
�nSû�(9�gQ㞲�{1n�)8F�H<�(gIֈ�������@$�g����Nx�Ac���v!L�f���v�J���w��_ �"W��r��h�!a����b,����G�(��;X���U��vZ9`)-G,q�C����׋���<�����~��o���To啕�i/�A�BVZV&x`�bJ%�P�I��#9�x�\�nX �W0���
F{?E��I��C�^�� �.R�f�qǬJ]:��xZ�@K0�����z��o�Э�2��|F�/Y�\v�+qR!6��J���S�
?݄�=3
nn8	�I׈-�,�����B�&��fl�׬L*��W;e9������x�_?Ҽ����7�����]-�:���S�����kV"Ei��R|�b���#�0<sJ�r���	o*v�A���=r�����o���)�5K4laN��t���������y*m�2�|4F�ݸ�U�؍MK��2&?3�&n�z�P
��
�?q�]FB���o���'t"B�{L��V��h0.���׉i�u��F*Ovy��թ�gπ����G ��L���)��B�蟲XA�l� �H0�kU,D�d,=Їx�y`�d�tF���p��
�����rGp����	f'Z@����]|�ǎ�Pw�63_Fd�f�����`%d��T�e��f	�"6�U�@���FRڿ�F>�e�_I(��k� ����0��!h��h+)e�g�uF7��reZ^�����6��'�i?��Q��Lt:����&L�iʠ�#�>7�\�|��G��GW*4�	onZw��"��4�����U����h�B`���
�a����c���ҷT�8��E�
O����^�`��d��J/B��C�/Ϝͣ4�VO�K^�>;B��g�4j[�M�������������~b�I��	'4��8������RVf������z"j0b�6�%�T[�&(�y�x�/�������*�oE�?�%�3U��.$��~*�B/��`C(���)���������bB�b��!Aj]��r��
*���G��)�)�v�u2�S�Gǃ���y�ï%���۶jO�d�!ats/Kҋ��6g�@�h$7R5�j��H'g��w��֞Vy�D!3�ꉰ����yt�I'�����䂑���w�\��M(L��xC|Uv�����o�d�8��5�Aȱ�gN,�i�b�W�@=��q��ʋB���AJ��I8�d)��B{HF>�8��Q�3�a�ثl	��9�+t�nǻ�s5`H���
���F���fIPr��d�e.�&��Zw��|�͒���:��*���,���BӴ��e��(<�z��w;|R��ɣ�6l���f��Q�S
��ϑ��+�����"����?2	I�0(����xp+X�/���nEdpsJs�yk
Z��t N&����ǆ�Z1M1��/�|}J;���)��
�tY�[@��_�P�'IC#g�R}_L?l�F�K���՟eC~�~����ԓQ/	"+eݟDv��4�����tv(���{e��P��~�;����)�ua�<�}3!�<�A��{�Pv?.X;H�S�~]��
Q5�K5���L��7��*`�J��}�����qe�3��ľ��9�ɧ�!��_�RG)��#U���^�<ew���N6�yl��/Yi;>���v1g�b���,�E�y(V�f
=4��U�n�l���%�N�o���!ѯ-�y�3`8��_M~�����O��ݔk02P��տ�\>�ŏ��b�J�>�dCz���'���0�h���֤�|����%J�{YdsV���\�q:tBI�1�����UO+�Y6���@e�-`�Q�*{I_Y�H�I�"ޠo�cUb�r�\_�p�s@��=���!��q�-��~�p5,�ұ��AK!����M����I��x�LT�u��Y��@�Q._��%�.�n8����ypѺ��|�ښ�i	�'�7\����=�o,ҵ:#��I���o��խ|߃۪��@T(@@��;.��F�oN�܆�ح�u�@M*��a5eB�S$�������U^P㔠�cU��`��uz</��8��@p�����Ԑw�;T0�Si�<�yM�����b����uV��M�ˆ#2H����t�C�m9U�ʶQ@�������`�,=.�@,��.�\9��y������H�����,f�T���jI������B4%.E��.CT�6��u41b/��d݌�%�=�RX*h�9��(=�� �cm.�ؚ2��z���5�����0���_��i(b��w�<ys��G����^%�A�Yt<�0ٮD��s� ������/�9DP[鈦q��.���ꅆ�}=B�V�q�4:")c�]�ܒ[�1�a��E��)B�I2ʿ�]�p4Ps�p�0A��!Gl�m��6Aq>�v&6/��$��6��
 ��y��Q�4��ی�MQ��H2D\$�-z����kz{u������R���TO���r��v.W��k�|��6ȉ�N�;�X"P����{�7���qގ�)E�)�'����ftbs2�m�㷘�45�sO/���r��R�h����W����)�!P�
d'����({+äT
�e �.Ĩ��~Z�o;���t�Jض5 ~?]�40�ew���t��ú�^p���?��h�.n^K�R��5�k�tP�!8�J���s��9IP\HG�<#�cu�9��F���uP�%�G!dl�1ߕ�~�r�=v��8(������� ;�r� G6�ɤ<ྤ�"�����A%K�;J��������1lI1D������Ϸ|S����~���ª<��7z)���{g
���K=?�E���U����_�V�IK����$^�Ѩ܃�qc��s8�����L��}���9NվW�0H^1>�����,C�PJ�h�;��S�4c�c8մ�S `�.8��D���)�ˡ#�Qq]5��O��a���)h���w�2�}4��i�AH n9�E�"�����T��':���Ph�-F}\�լkr������olӑP��*|P�kK�G��]@�l.�NPG�{�G�h��S��
��%+���(�O��Nz����.���@G\";��N�:f#H����PS}��`B�;eo�k V����	�Q�	��}yV����52ց˵��]>�᠒|�&���¦F�Q5m�-���I�/f�7�����wX�m@�w���y������|�_�C��`�C����4J�{���X����/�f�ǚy96�t��&*B�Qy:�(h);7��NK)�9X�"i����"�Ή����gwdJ�����[�Pb�Ψ.�z��}L�Hd�iir$Xm#��!�d -�o�G$R�Ow�?�X��E����Q/b�.��Qj!M�	;�)	�ݯ]�S�f?�.�b�:��yӢ�ƚj����J�ۻ�8���p/�Oq$_:�3rNmψ�F����|%�%��I�xZ!�"�c�s%�`��0J�H�	{ƫ-��?ɿ<�DSEXtt��غt�U����~�0&*L��)��@:�YQY�]jYI���8k#��J��>7�\�޽��Y��VLn+a�%�`�u6�2<���e(���Â�4_^�Fp��斕����&�����;�[)�Yx���V��\��r��o��֗i���#(�	k��>����ׯ�P1�3�'�8N�[�ir<]�U��F��B��{f*_�~�~i�q����u?I�9'��G4E����ma�@�f$�K���� �,��&��iN�%H>�A�搲�}����-|i���0���,1f���$���N�ِ���6����6+�z4t砾Z� ���M��e���'�$�v�� *Wn�W����z�k��,C��՚	Y>,�R�T�������_i�aC8����o��p�����	)X�r�Y׼S�Ĉ��y�q�^J�4�ke��E��	M��W=&�q���Z׫�~�H<��0dϹ��o�<|h/,<[Fx���-�ʇ�͊��8GO���0|L����}M[�Z��t��<���n<hC�̦�w#�Ճ����h6*���X���W� L~qփ���:�����U��C.b�
;�Z
t�.Vw�3��$��䫙a�}���k<Pp��P9����z��lh��i�!}d��0'�'�����(!cV��x�D�o@�i�m�R;5G����)�ɦpu������)#���4�2S��(O�H�B�)�x~�Ѵ��5�d�e����c�� ���@t��Ĭ���B�����6%�&˩K�TM]�ܑ�_��̈S���� ��w .�����ޤ�Ŷ����}=s�c�����|���t��E��gZm������}3�|�ŏ�w3�g���(�tH�r�~��YL�tV��pr�>�<U~I��"�������t_��hK����rL��=����1���!p��D#���Sv+�#��b;�U��H�ݍ��/�q�iД(1��֏�Bcfv�XV7
B*�厈��L��4�ʓ����8��w�s�Fz��Rp�6�&�ˉ��k��?��7�h�cU��V �TK&/!�������>�
m�/�!�(���M�y�:��M_� �%������z��Q�
,}ٛ��VO�X"U���:#�˃�C;����ٰ�7��<�ڹ��ɓT���y-��{eǱ�E�?Ex�k� ��<V�pN`6#� ׉���LM@5�%�CJ)�3�]��Ua���z�ky�[���'?S�'J�?9�� ՘�f�u�j�mq(sS=��X���]����j³�?����9�p��֡,�����61h0`�F 	���5�+��: �DF�B�&��d�Fm���6ӱ.d�܍�;�4R@�H ���:o��֢���N���8��/����x�oϟ���z�h�i�L��Gu9d#E���K��<i�Yd�r��u�A����6�p�J��>�ޯ��^P4����wTfk�q"d�9���]�2���BB1�]g��3S�ʖ0Q��F����}:�I�����V��A\�d�㥤�G3����}J%��x�P����J�Wvmb�5������J=h�d!"��G�r�}� E�߳�U$�^8��bkt(� �r�{߱���払��a��aa]�J�u����N�TƮć����	���&�>/���6���H''�x�M�:A\e��������	!H>�O�,����Y_�|{Z��!P<0��&�6"0�!���e�z_b�#>e{������������� �C���Z)d�"�ֆ\y�y�S�m�
?�Ax7��ͬԨ��0�޹S]�9��������W����l*ַ܏��:�²@=կ�]ؓ�̳�O`�I�ֻ�%�i]],d)�P�_5�D;��$�}�����(�חEo�驎�0o�8�^/XϨ��"�:.y?��m�q`��iP�2�Z����P<�� 5d�j�V��h�WK��E����[�� ��3ş���V7Q��%����x��u�W���9���n�n(���yO)X8�+�]��߇'j��δ�B�ĺ�G�r�g�	qEʭYp�������7�. }����?�8��r��{��V��\F���;Wa?�2[11�S�r]Ն1�WkŸ�B}<��+��y������@_�JM��o�	�'VJ�z,�2��qv����0�~�dy�	��hQ���rM�-�Zp��#��t6�����R�
�P���
�l����,\JĘhzNWeX�'a ����37�@ě��"���u��8�8f�k�ȯt븿^�wN�5��>�M#�h�/¶�Ё����lD��s�A��_�oIg����K�|C#�u������:Ԣ5�J3�uy{�p�Q�t�X �GY�퍫��qY8�|�S����E���K�K1�d�������r�E�l�ϵ���)�%��d8��AB1��w	�x�B��=(/�	V,�A��}m����6~A 7Ϭ���gt	��HsA]se����*��V$��S��G��������0ė�rj�Հ�����+��q����	x�A��Y$Y�]���ن�u˳�� �Cn�p�"�ԯy�W{G �#�a���u�&��{����F����s���Z�j�Myڦ��b����t���q/r�6�-���$h�:�n�Ȓ��	g�L�����7���j��[(��[,��i�P�}��J��[Y�84�皲�*���mw�|��|��&aq��7P,Ǟ��.9Q��q/a���C�������}<�!�ͱ�b��JP�]��%i�U�o�F}��=8u��Dk��%��T=kr�GYO���˶�T��f}��|��e�f�c������7J)#�K�n��C�?%�����6��|��P=�8�\jtAj"���c{]�Eᩍ�v�����"^�7Af|�de%���ȹߌM��|�?�G	��CiF�$�`�	 ���o�����k^M���i�z��NR7ŝ�a}��Խv�� 9�GJIU�=5��G�"��G�!����Pը��.ZDg2�����ǧ�o�C~K��v�L�F�3W�Z�ϫ���ԛ��@�)�Z��[g �R,a�k�`Y��H�k�0���D6v��(��P%�f�"����S�'F�*�<�}ȥՕu	6��1��gv?F��B�Wi���R�@lx���Ҙ\��/�����i����/�B-O��l�X[9��мbUv_h�4�ov��}G�Vf�����AN��FX�t~��6?�2, �t��!���f�W��~�����>��������4�)�M���H/��ʅ�G)����na��a����Ox���q�Q��GDEoĪ�-��8����r���dfP��&%���s!ex���G`I AN���Lt/)�2V.����<���l����a�!x���3;��Z#��3�u"W�$	�@{�@�h�A��7;�� �K3�G�`��$t��d`w5�p��%#�+�P�<�pC��� `��M�8~9$~˟�Y�������7��P��ʊ:v{`{��Lܑ;�UnY+٢�iK���o� >V���� �O�rXadש� ��0�XL9A06����.@A�]7��PRM��1v�'ށz�X�y9�\���ԃ�sc�а�@���1�ȉ�A���z
��v4�/:<�!=�P�� ��іYV�̲�	|��n�D���G^U��q�-n^�ŵL�z>O��b�E�8=|ض����,�
jr�������O���Z��{�/U5�B5,h|U|�������'3�b�2"</֊�(�(�'��!��G~�)S�=�*�ipR��:Cz�A��y�(�ŭ�,k?ԶZ������֌Ss
RġF>�PG\9
 �b1�����G��[N1�����GAN�W�����+��̣)�i�״�+/����c-�-�@TK�Ajr|�Z�����+�~�F	 ���*��W��5������׼?M4��?M���u����:��}� Dֹ¨���M���XmU��:a-W�k���0�|���oZs�GD-� ��D��U��-}� ��?H���0����ܿ�G��ͳ�q��bG���}�@����6�)WƸ�w\�ӫ4P
���޿k���k�]q>� ����{�`��Ot/#i��qr��b��~��jr�yvd�<l�����ᇯe�V�AI>�w�4�0����^�`��v�`��S3��Q?�<��%~����V�!iۡI�Z:#b��it����e	`�Xw��cY�j�،ʮJH�:�җB��	���+.�M�P��J�eT�+�{;e�%�X�B������bk3�<A�"#������z�cG`jӒ-fD�kv�2�71 n� �R���hOpѧۗL�Ie�b��2��U*�C�]��S���QJ�q�m��`;�W�h�v�:p����7��s������AlƗ�
�ho_�@��c�e��N-8��ACT�@TD�����Ӭ��Zn;A�6 ��Ԯ)�9��┠T|�����QmY�s�o��Uޣ�X�})yGX/{<+�uiD97��YH�y�Z��z=e���{}�v�	C{��^
�s�[z�t8�0�c�<��A���0j�Ɣ��������_�43��q�t�iſu;���z�*��iH��>�A�%0���r�w#
H���gs�
�C��Ր���:�x�����L(x�@������9�Xvر!ݢy�sq�}�-X~>�+;�1��r�P!Bp���^}#JeK�K�ndX�z����˘�y(w����I���5ld	�F�8��y*�	s�=����^�m�A�'�+����f�W�
F����@]�CT�H٤Ŧ��jy��H�A����m�g 2�<�c�.3�G�k���0x&��r��f��,��[����f�o�X�[H �0�{�M����L�@Lʼ`�}��[yc���n+MM���ʩ��u9*�*1?T�
�+�Y�B���c��P�aH}x��C\4FP.��� lV� �#��i����剨Y�\��tV�mO�e.���JN�����j���m?�L�����|S:�(3Ȅ�]��~7ھϕ�I�~���|�D�$<3��s^�-��\يXe�p�������@�&=�8�Y�ި=�?�ų�'t��D*�9z�Ä�T#f��o�M���H��zH��D�l��~ڲp�yT�<���ܩ�)��M�����%���������bО7	/���AR��];�fL,RZ�'ne\@ٵJ"W�<~*�Z�9���̩<� z�^�9��G�S��leoTŶpu4��o�R.�q5p����(���0y�������z�	���Pm���T3ԍE{r3��<�N�t������R��_Z���z7���s�h��ۀ�*0�7�$n�ľ�����.{fV*.b�Տ���唞��v�k@<M����t�����g
d��O|e��i����[J�Q۳�Pv�#�������fq�뚤��]޺7;���!�u%Ȃ�&��:~���JS�.מXy�g��
�&?K�N���B��ɹ7d`��?S佶�J��nd�d���]yB����R�;8�����M���?�a�.�e�	�x�~䚆�3?o �x�j�����V֪+3�c����GxFmF㮒�$���k�<�1��,��[:�f�#���!�;�
+��[&�5�5,%�o���9���	�"�Gv�I��ü�l��ڱ*���w��A���?Z�T_�'�$`�	c��&�@���:5{��Y��ʄ^�<��\���i�S��6�$�,^�a3�sxs�}*c�,�b���n��_|0/Y����T�\��Y���Sf����#z�i��M�s3-�{�})Z?#6�٩!��<d~[�$�>���n��.�s}]c���ո�{π�zg�t�4��^�'E�K��v�L.��p�y��Uvӧ4�����6J�jw �q��c����ݤV9�T�������=����		��b��B�tտ��2��"�u	ms�Ѓ7o)�"~�����4<e���ݵB:墼�t<R�a��R��$��s7M<7]薢ϟy�?c'ߋ(SW���wCP�fO�,�������^ԥ|�my�����Q�Y<�<��Pw?��kpXD�El��N'�b��B�7�:c�U4���; K��d�hV�{j =�İLa�O.��}���$ۍ�Lv%�G	fA#�/���7c���ww^��*��X�E���TV�����
�o�~�8��~�Hc�f��Lp?2�e&�H?E�h,��R?���U<��X��������PN�.%%��s�2�.���}ad�_��-���ި	M��X>g�N8�cyQ\�-9`<��272$�4�Eux'��]3�x�E���:.}�Q����u���q�䓡n��Y ��PH��"������c���yQH�m���ڟ��ư��B��A���d�s?-[� ��
O�p�T�Z#�ʫ�
��b5�Ω?13��񷖁�����1��5���҉����2�x#Sh�7حL$��iDj�L>�≱O�]�y�����b^N��Xȏ;[ԖK�j����5�<���qi���D�t��ӻ��%H1�E�c�&��𜹘���I%���q���ˍ;��w��z�:q�:� �;�ږ�̥}D'\z]r���kn(�n(u=�
�,8����f|���6L�V �-�9%C�΂J�.���2$�;r#�N@�/�?�.�<�x]�;,;h����-�XsE����흷*
?�/2q)O�@

��qpo�<Pb�J��jjK�%��eA
��>��im��P�h)Vvज8�,���}���"�_�4�Z�Z���g@
ҟN,�$p���C�D�
0'�.�N��u
kC�<\��W���x�]�6��C���/��
�K20���h��=1[�jN�#�-�.�r��'N&Ƃt�̉P�w�;`	޼>�#��cT�~�7\��:�s5"�u�8�R�}�T�&�e���Bf�4���c���h�q���ڧ�UW�h=t�;1F����X��w�H�b>�8���y�?'��!��5'=ۢw2������uOa�|���N�&`�hS+�1k� �=B֢mG��T�ޗp#;,�ʵ��s΃��ʽɟ7e����i� �/�#K
-U|�5�1(TQ]@vm}��&(��W'c�(H�S_HH�}֪���Iǹ@
�Q��鞽�{i����ϐ~q�t�
>W�ؙr��6U�X�1L�t�*�yN(C��Ԣ�	\�bxi��P�rD�&IעDR\k��#��-Gm���G�2b;����.�.g��I ��C>�-��?������h�~�;"�໇-�>H伹��;w���cA-�ð�i7�Ɓ޽	r�k�A'�-ea,!��֕@���ut��K�U+���10���y�fߧۉ�Lrn�c��2��;<������~�
p!���f�-r���)`Av�)H���F�+=|D9���	�ߵ����^�7�m�2��2�@g��5�y.��-�����} �́f�rg����S0���;�ȫ�&f��� N����@w��s�ߖ�V�b" UôK6^��Iy�������M���h#-�栿<�&w��1����o�T�T�ӥ�� �$Z�fH�޵�^����:��\�R'�G�	95�Hm�_��ÖuY���?����d�b}�q$'��U���;-�--�X��`��(kt[�9�7�a�u�����ljV'b2�\��&!/Q�&l{=�=&��A��e����s~�I]��	jLt���;h��l�a6�ͼ���-RbD���gֈ�s��"��hé�H3��2�d{>�������FH	^}�vR�[�ٻ�\Y��}_\��{��GMd�d= ��H})6Z@Y.���}�%�-���/Z��eQ܎��8�����1��#i�*Q�E|�ذI�����,9�G���#rDH��nbZb���e�]��8�F�{6D7��}��BIr�}d�Sj@9�N�6(�6�#ʓƻB��&V2.ivi�ޮuD�<݈�"����Emq��/��;S&u}�E���4��5OS]�UF�9n�}, ɕ�]L��w���"�f^����ʹ�)oѳ��y
��0��5FY����D�A;Ӯv	�&��ļp�Tg��,{��Hj�N@���3qjxR��{�]��ȑH�O�~�Ýsw���Mh�^���/�)�f|6�E#�J�+T��m�d��+����٨x�Ј�B��W�����TtDO�0**�7�Ү/�2f�_��Ox[e����0��E��l|�v���s�`��H��ƛY�����IB��c`Տ@�Չ���.�@${��p�g9\FZ&�P?�Yȵ6J��"����>Q,�:�GZ���N[r=2(�-{�u�UX��2*�X�7h*�T����u�ڰ�amޤ���U����A���I
�QS?{n�{��H��3���z��ݙ�A�[�M��l����ǥ���Q�����	a�V:���h/VO�V����n�ɞ7��d��D�p
N�ō��	�h�m���S�H���.z�u ����P��Jxg�w�I���J/�v����xg,�.qO��� \47�g�z�E�hqpE{�S�u�2c���6�޻ѷ��3���[\g��h{�/�;3Y������xѾ�y�U+|�I���b��'q�3��
.~�X�`����e%W��vaU�	) ���2O��{�e2��eP�H�50C��EU���x(}����Dݱ�޾��<2�6�P�ϫT�&���>���9�k�q�A�ms��^�c�C#ɓJ�CL׾g���L�~S���<ƼU��B^9vZW�D	8�6)�E��.B"���w	��BQ�*o���}�-��^t<K�ձ�!+���6�6���<z'q��+�A�����5w(-��T�&|C+��Ab��7���\E�hxS�Nߥ(��N���}K��d�Z��nM��6bz�+.����}0,�����_鰠2	�d��m��r���)[en߇ZȾ�� �pPL�%U�ψW�
0�e9���E4!~����IfjD@�h��7������c�B1> �����RC/@��=[B��g��3���h�!*ص�� ������]�70´2-�w�V�;�	w��@6k}퀣��/�-2�ݞ��'�>m��B���>S�SN^����������e��*�G�N���tIQ�?3�������}�nʭ�G,��e�2ȷ��BR��P�,���m�+�#-��ڹ��х��. �B��ԕ�9ҸF��,�����W:�̯��H�,HDVC��d?X�����"�e:�D���ƛ�=��_����{�q���I>�Ͽ��]{R�� h$�p47��a�PəJZ�M��CN6��*�.�ʽ��O.���}W�D�9f�m���1��1 �N&~���]�:QzǕ~vLݫ��J2|�J��L߆�?��΋V��("��$�sdM/�D��[tZ�A�^MI���ֶl��7�=XN���%�M�l�T��G���x��4Pr�paPJ�j]i,T�W����5��s�A%LZ,�b@lI�H�D�9�X������YrĻx?����[���o%�酧iK�>����$ 㵠�h�C�=��	��s�S��u&���
m��i�4���v��:���T����`J��k��S'J���_ԞQ�#����ė��F8��* f�{��NjxFt���Fid�ӝ-���g1,�	R�M��$bIZp�Ih���Y�y�םV��9��j�=�׃�* N������\q��,���!�c�6L�Y�Vv�p��mU_r���BJ�UV��Z�� ����d�d�資%p��b�x�P5�o?62����e��V���/���<r �AGV��;R#j���c��7�(���,�1?*�q����I�{�x��B�
J��YI�-u�-W�y����tIX�ݫ�ͫ3Gv���pw����X;� ��]wWEYĩxP)w���I�:?�ޱe�x��w���k f�{��%"�6Fe����P6����u� U��h�+�gC#a��$u���Iװ�]��+.p�L��3M���f�x�}�4�E��]�E���/Y��u /t���rٽ��g@lhl�ps�KZW�	��k� �M=5�P ������9���1�.L5aI��4{�>;%�[4!�����k[[d�R�7sb���;��II���?�Ϙ���^sX�}��4�&��eFrr$�A�I���`�4�c��m՝�L�|��󪦕��W�
����0���EXƮ�ο���~g	�t��s�jL2����wW˅���Z���=��6��b� e�u��a���p\���IAWX����ޕ 4�妝���C\�0�RA�������}3t9��ɔ�!���`��-CB�)0��+���ǎ�S
��~���Yp�Pu��ˁ	��1R���#np(���&7�=�{�D�9�C=�l���)�(YVd@��*/���:�,�F����0Յg��ɋ�?��|�CP��r6��Q�U7�����[��^�
7j��xPU>y�r��f�c�ď}: N�KX1�Br	������J�븭`���`�6$G�;�L&��W~[�b��=��"�kn�d���$��=�vH���s�Z�ŁW��Hz{L�Q��S��zs"?�j��8kzE��[�!2��Y����P�Qux-���b4!�B*oөlg�w�����ĭ�Lt�x;	�)���M�j�i�(\����t�aG��8�mG�33rN��E}@��+fav�J�r
�- �E���0�a��I��O1��<�K&T�E�a��yf�C�9'��S��XV ������א�B}�<��~�U����1�ŷo>�waUu��?$Vy�h=���ץE��8C�k.1���C��W�M.9���߈�>t�tm3�#p?19�����S�ژ-��F<7iw��&J�`Jqõ��a��?�œ������25>��8&�vX�>W��L%H�j��+���$�������e+H�yǪo!_W�C�b��V |�Q��*��ֲ��[�jVFc�%�&6��lv�ہ��;Jv�
bgi)<o�̫侶� ���;0����d�ɳS�Y~����8B��_�����>mt���B��S;��Q��$��Z��9���H6�$��`��MFf����Xi�I�!�k��>�0M���!
<3�=�2M��!���.�8u_9�#�*�9�� ��H?_�"5��#�e���t(�����U-ۈ�I�p�!���{�~��N�M���]er%�!N~��L'�wT�	����-U�Ǣ*"�SҒYy�?:T�)|�3���2H��<��t��u�s]��P�sr*C�v
�ښ�4�T�()*�Z0Sp=���k:pi*�#a�bNJ�[ͯ�J��:�����D ?V��*��B�&e=�yI��d�G+����U�G�.7�(��|���)��E��Xc�ʷ'�n�<�K�Kb�U���AB,�I���D���s�v�m��\��>b'�	�F7�0�ܛF\[�5�1>Hr�����:J18
<|}O�;�i�8rgv#v���}$�H*D�@;����W��V<�7�%%�WN��D�E�If'G�N>>[s��'�A&�W\�J'�a�iNq�g���}����� �ҩYtY�u�x������q���}��-����;�V�O-Sw��$LS�%Z?o�0�1ȯvLͫ�'������?�+�cmڳ+�/4��2�$��G'j����b~�d�o�Be\K7<��.Bh����e�C>~%{Q�k�}��h���sz��c�m�N�H���̀��܊�$� �3	�=W�џ2p�lqG�C�I���U1�߻Q��3���"jFmZ��
�'�v��-��Ww5��WmҖ��`?R��~b���8%3d/)�;^�� ����D�y�l8�,���^=@�@ѷ��z�~��I6o�~B�ݔ'�ҏS��&�ڣR�Z�D2���(!P�{��f��S'�n��Z{���';��Z��/l�Ώg�	��Vc�+����u�	:h�"��6�(�#�j��p7���0����9Ys�9���M���� �%��v������6�� ���%�$E6�ŷ*\�nI��"�B����+���K��t��R^��oZ�ά{�ZH[]h4)㷺-�z͖��0����45/��[3)y�^��UWp��([��pwA�_%�r��wP�ym�A�^�F���fb���6�����~�%������?�E'[�Z|��#�-�=<�I㘛Ba�"����}��C{|�����<��z*Z&!y�k��3�-��)C \)���x�h�q�3���y���Ʀ�^֡=j�I���Jʝ���h��x�*��,?� 1+~
L�#�SB�-Ǵ�R�������m6  (�
��DM%	!)%Ct���e !���Y�/�f׭P��f���+>i��=�2�>Z��Hړdc���f�{k�5�%EP(���H�#��<������Cq��������d�����=����gn��\���z�R�I�����6�B�$^��vӐ��~Nf�nj���4j�-Qt�(MϖG���D��QdTУ����8��p���t�x�Q���V��O�I�t�CIa7Lఋ\�ٛn�=�;�:`�nZ1��p���DGb�Y?uF��*�?�w׉�>/�E���8���ġ�Ȃ7�~M`�p4K�����"zܗm���lX?ǇE��,�l��yܓ��I����2�|Z6�?��:��!��?�6x۩����H���#�"ũ�<󶗗�-��U��R7�GUC�<���?���m����C������]��_/�V��/Q����@e*A��?���o�ax�� �3������F]���y;N��[7�vƝS"� v
�_����^�3��.B椵�������1\Fǆ��w6�MZ�"^���G�sq�؇��$�f��m��>�ϚS���K�kw�5�p���t�[ErՈ��: #E���:�EB��)_h*hl�7'��@�m�踁�Y�v�C��(�`�ʔ$�g����:���_hG��3�o���DEL���&흈I�#j�ǫj#� �XOY�Yg>�4᭞گ�^��]K��C��P��������'��CؑWa�bt�K��5��m��1逷�1�!�2�38�"�Jb��@��J�ε�E��7�(
��&Z�����-��C�>��c
��� ��5�u����|>������<�!�}�?3Fy8�'C#�������M�\�ㄽB�����O������n.<��6�:�@e)���Ƴ}��q
?�,���Ø+�感}��~n*m)�S��oKb�����&��dkؼQd�'<��5_~a��[A0����{�����NH���ާ<��l��a�~���p9�u^�R�l>�\���g����@a?��i� 9V���!��Z�&�?r����-E�����w��:�V2fcødʇ��Fzc<}�건IrP_�r"��ʱԨ��D����'��������k���� ?��b<��*Jyz��!E9�꭬�X�����>9dO���}Ps����
��֝q]���\�<5O���9K�#���t�?|�9R�J9V�!�?����n�Σ�j�cX���2�����O\�]R�޺����g)��������|O�f#ϱg�QZ|46o�V�N���5�R�k��%QVMV��禔rg��E�l��ɀ�ѽ#&�X�͜�I'cШW�� ��T�̢�&��2�^��}�3��]�Ȱ�j+g����+��\Ͼ�C֢)h)B��a�a� 0+�����U7Cz)�C[�8
y&#�V%qM L�h�O�n\M��h�I����w���u�}�'�p�-��-Ҳ��/�Wa����Y3
y!����bnG�C0H��J]�k�P�h:��<pPl3�b�ƭ�t�F��)�4��.��J��H��t6j�F�y+T�e�a6�$�מЃk$�"M�v�hl���
A+�CM�`/^FB��Ari2�kR�ó0]@�=�����/�d�fe4:����$��t]��	�
��ue |/1x�T7v�7�j1�rV�Y�)e$4 �h[�ny������y(0���)��������J[1V�G��j)����Ur�����(i�޿���7�����
��Mry����e^n)Ҵa���@���.3�:}���� 1))W
���;�[_��`�@4��t���sl�ѣ�ׁ	�K�\��
C�"�&�PI	\���_ ��*�ݭnѪc�l8��o�w�t.Mءa�%�Cۚ��E�8���T�P�9�1���x���*P2B�KK�4cn���i-��j��^� W�:�㩊��۩��Ӥ�������Pp�vn���XZ�5��3��"X�%D�W靿7h�e�ى����0<~U08~.>V��I������=�_���T��JР�E��ԜTi{�2� �Ӹ�����o���qj��b�Ҟ5t�
~�Y�����x5�i�i�VVs��DG�L+����-�5y\h9�ԛTQ�IM8���Ա�,7y��lL�_�(D�z��g��(�
�;H��,o[�s���UV:�KU�mGp�%W+(�i37S���F1�!�.�D,\�S��*951� �����^���ī�1`��*λ\O����T:F�h����}��
����L�NZ�S3��|�W��s�1�6�LI�l�7��α73lo�� m�cod�$�D���d����]n`#$jٓ�:ABQM�p|�/5��-9���Б/q7��	5�5���R�%�W��h��z<4Y[��&d𹙙��kV�[sBޡa�i�9$ğ��6���a�=�vh����+Ģ��N��M�?5���d����v�ϱ˳+�uם����2;��!��ɼ���N�[�j�%^ʯ}(y"�����0�A�n����˵��r�$o:g�hf_��F�l�Wx�O���%�f	
V�Q�*ѵ�j�w���W�U��p��G�߸y������V����Lj ������$"�c{�{��u<Ojj��䍽v7�9&���->,��AD��T����\������Dk�����t����s2!n��F\�ߞ̭&�6������W1���F�а�� ���.�!5d�ڸ͓O������z���x�MFe���[iY%kH`�z�,���!�2�TN댃nw�%r�^<�5�k�3>Ny�ν���%~ڟ��{���hSm}���Y��ёڤ�:�lȆ)>R��,Q|-��F
ګ"%Uʀ��M<	�9X���4�Tu+� �2���*�v�M�9wI��U,Y�&�<4{ނ�`��L��㙢���[��)E��-y���$�	J��ܵ���*�:38G�T��;	
��������V�C�Ԩ"��Hn���09�r�4��IJ����#�8�)���e=���x��L�����/!a1N��k�'�洮:�'��ab�do�)�9�8
���}_�����y��u���;�����]V��	R�*������,<�y��=�\[����?p��Xd���]J4t;��L��u^�
��+��w��%�`D�K�&�w{3�"��+���@i������/J�t�FX�b��8^�Q��.��	�4Ã��+9�v�j�3Xu� l-��'�UeȮ
ϩa�^�x\\�Z��8�@S���Ӆ^\�;r>@�����3��ԙ/Ӓ���+~r�P	���8�0
�\�w-l��~vc
e�ϊ�d���f��o�Ml�5�(Z������d,֗@n��N����^���D�cW���v}hu�Q.q�}���O�6�&��K��I$L���fߗ�����b����\�v'�I<b���S�li����6�E���f�߁�ZU���.��`�>W�0"��j���:���H���~�XY����>h{�mao�+:��b�h�{��^H7�����Y	5zm�!��H�ά����j��ڨ�W^c/j�5�� �����h���م?�H�k)>����//����@���	�jo�[.����s�wyW�����ԧ�_��(.�I-D�Y#S{?@/�VJs=�e��P6K�Z���Z�f���؛č�ʱЬ)�z�"jf�8�!�$�5�?��墀3���ԀшD���p4��胩�%$C4+^�z�|r��Ě(.����Kk��s6A?Xꖐ��Uu~S�/s���6��p��y���[�2�U>	�Wp�]�؎�BHF5��z��n��:蟏M�$t��cJK�Ţ�Emh@(�
H?�`_,[��]2��Y우
��v'�ή����"���=HcF�c�G�h�����j��N�X(��t�f�b̼A?��	���t�4����!ɵ��=����&�ǋsF=�h�do�8������~��N�;,���ʧx*
��� !�d�rJ�M������H��$���^��C���ܙ.�����V�5�WP޽�!��<�>���~�6���q��� 
Z.�k�=a�����C��G(̱L�02/f��Y�o�$�����QJ��~�P(�޿�#?6qda�T+�3֗��rF�g3�'���ǎ|ѻצ��Lp��:�����-/峡�:^N3/���q}�]�d�]��#�+�e�:�s�"�N5��s����I�QM����z�ܦʀ	�%��<&��h�sm�D(����21#u�IʒM������I0�������GߨU���é��Y�/)?{�����w>�S��@{��X�$c.��R��w��_w����b;bB<N��\�8Nf8��-��;��� ��29x$�H|,i��al(����p�t�w���贃��,g��5���=�����ۙN���A�����sm=x���'o���Y�DMb��o��!�m�vݐc8p3��1wF�܁ݷ3QhcE�P9qD�3aB�p$��z�W1��]Q�*jocf��w,`����f�XQ4��~�j!lT)VQ.gY�텃��Ɲ�J�TH�b@b�t�㛳�����-	s�Za������RXV[�:~v���?��)���y��o`�nފ��gΗR�F�T6��˛�&7M� ���m�tJ�\I&��n}���/0���?�] �œ��nW(�3�s���� �ߴX ��b�v[cBǆ���x.��]�(�����m�Y�6�Y�����������L0���|}�rW\��Ŝ7�8���|����_�,y��Ǖ
yR���BW��q�SO}��ƞ���
�7�����k��6��w8�%J_a"�^7�v	`�q�|m��w���9N��a�>0��c�ꑫ�1YT�L��p�[,1���J����+��6��S��;�;d���9&�S��Wc��'�Ԙ��G''�'���&V�͜d�z���Q���p�}�{�H�g�8�`5���H���۽�7W���ט��l{�=��߈�1�<`�H؋��8ZJ2j����"��(�p� ��q2ߙ��(u��uB����85*�(�)��ą���s��W�*^���P7��!]g��Q���/ћ�a�����ۆ� �#��;Q��
�x3>{h���%]�Jm��,NeQY�T�C�m���Ս�N�6U/�<�] =��]E����P��y,�5b_��{-����t٘"�Q�@��C10�@w�
]�3
1i�h�K��V8�k'(r��ꋝ���_; �k��u��v�MJ*H�`O�t���Y�Ƶl_���H^���ٿ�@����E��4��qT
��dz{��@%�E�[�p�	��h��Jw~
~J�a
6����*��
�D.>�"�"*(�&�E��?[���m{�������y�f쀉CY��� �\��x�!'��(��#���Cd5�)"��7o~XttX������r�}%�$:1W��k�����9���!')��-�ٶ�.����	�h�8A���@c�N�.,�$�Mِ��|L�=���߬*�j��� ��7�R��7 ���(p�2�+W����(tׅ��� �t^:�F3xȱ|�50�H�j��mnh5�>0.y�>I�6c���uo���ܥq�o�X����$���y�Nx�6m��T�Jl៽���Jb9�*(�� ���E�c��5��r�O�0�Ė Q��F��5ۚV��{	���=��n�t%s��ŭMZ"ẞϲ.���_�B�Í��$� 2=�G�$`��y|��% w.�G9��jVi�V�t3d|�� ��PM�.�����:�߃_r*P�Td��QM�@.(/>�BLO�<������]nQ�[��_��RڼU�P#UD��m��	D�M��~��$`�I���)J�PL՜N���N��tANY�r�\5�K�K�������W�?����r�!٭��#�����ʼ�,s�#������D�u�����aم7�&a���]�d|����v,^5S�%	'$�K7��"{��_#�k��g�� 1�O2��_c��$�A�!е&��{���R�r�o�3�w6�U?�Ⱥ�8�ߟ�{�k(�݂���b���9�`��@�â�n$��!��t~_U=�Z��-����mm�uAL�M�������P�'g���0��RFy���I�ʼd%���{tG� ����x�Ff�o�Ո�e<�9��}�@@�����@�މr�{�Fc
+� ���D�&�邐��@�,��]#j�9�����T���k�V�/ֹ��!bF�����B�P&�+���6p�1� �D�lw�h�@�x��ۚk;nrus<���M_���+o�t��WMJ�ʴ���q�C�����$B� ���%�Du�����1��e�@�#>��(��؍҄e�����Dx��r�7Q�����m|�/X(���j�����wb 92��{��y%l���w�OW�R�{@[Ф�	�H��L�O_5B+ښ�M�7��)K�r��N}��}�\5� ����.�b09�Ԃ�gCcε�6F6���z0������[��?�@{�&w#�j��.Q#g	*��i�M�#$b'�>@��c2Gz�lχ��|�z���Q��0�q���j��]�K���'��#�aH��i�E3Y
���oW?��p���uL��-H"��B�<Yt�7��[}������-^V�NMv|��4_cM*}�(FH)x�gs,�W��|�}P0o�3Ä3����k+e��nTjк.��x<
��)�A�pr�r����ۜ��#6��W0�r¨C���hv�%��ڻt4�e>�J�����$B��a}<��������!�ĐmJ��ʏe�zhŤ0�6�u/u�����b��s��mp�a�
±�ߘ�/�����~`T��7�[6gS�y�8���.{��>���a���n�QBV\!�$�:L/���=��y`���f�/T��/�b��%/�Sdp��B	t��d8F	���\C��ɕ<�,�x>�[��&)��JC�:A`m��v��	е�d�zI��\������_�,
�k��ט�L�K�����P��9B�o���':��%���e��̛�S�>3��}�a&e�*��G����Ec�z�жф�Te�P춲ʢ���l�SL�#m���M�=����`�zS���6��[�E�(�y"�%Uo��\
p�"��C��A@ڒ�X�� ���ӥ��� SؼӚ#��+A'�6� �C9K5(aK���$!���T@x���6*�����0��ӓ����\��m~���\	�bn-���^��dm4��:F��ۗ�p���.m)������#uhX�I	��"�������k�@�ѫ%�z��"ɋmA|i������{�"��6�������T���%�	.s�yCKM������~5"��j����J���$���� N��u�{`l��/�~�8i�w��m�c�H�RdMk�8f(Z�5�w���B�c,?ժ��ܭ��@a����c�?x�-��[@�xԒ�.��z�6o�vSfM�O/ᎅ!���"F=�Cq�4S�wu�~�?y� ���Bv��f_F{���&+�cf3(Є��A��?=/Ir|����ug�1
�*$rB$��=��X�����m��n����:"��u�*����a�8+H_t� �`��.� 9��v��
p&�J���(���r�	Q�A�A�.����~ښ���D��$P�4�<A,�(�"`�'�F�X �|A
P�N����|-�������st��J�[\��3}���a�8U��U� c�������OX-5H��fr�H��{R���}2����#cG�� Q@�ލ��C ��2!?6�3�q4��C�	��>�,U#�]7���T�@�T6�&��Էu���2<,d����I�1��h�FӰ�<� ��V�"��������K�fS�熟Ё���|P~�� �$���W��K�5��#I�Q֫� d�
bv�FBT���,�\d��8�|�D����34ҕ!nL��S��A���x���*�J���|��^2�"��F�#M��øL�!���O�O1V
v�c*�xs@�r�bd�z�T.���g���io#л�eY�Ƣ&���xu���6u?�5���E�����{��e�-?]�U�١���v<�@	�Փ��H&����.ެ��>5���*�@��h:%��l/��u��w�YE��#x�3&��`v��t��غ2����i��yHb�Ed����\SY<Y���48�O�R8���>`��.��ܧ*����[)�J+�f��ꥪ.�[���E׉�"�
_J�UCeL{Ɵ���2n��Ƃh��(U��'lF񄿒Ϗzb����``�?��Q�A�C��O�k �*.�����C= �}��UK[�,�j�n�`t�N��Ȫ�G����c�ϟH[��}�*��	C��?/Yu^a7���͂~�w�;$���uȗ�(Kio��K�5�$�a�km��m`� ��*;�IPA��j��c6�q*K��cS{���<^÷
 ʜ���c`KѫA:Į��w�T�B̄Y]7�|�F���:����jrX��?S�5�1'1����M��u��@gvM��|,�f����U֍��}���<}B9"�����t�ӈ�+hԑ�z�Z� ˌ�<�v�H����(��O�Zsx'���~�*���1��!�F[H�h�ƾp��(q,뱩g��7�����(iN��|�1A�Ӳ�Fɚ�� +Kj$5,���s��F/-n�ԉ+�\�J��>�n�gaaEn/����9'�B��sc4������=��	�߬-�|�2k��������-5v�V���E��X�ҳ���_uǇNZm Bg�S�Ƹ����GU"sWK�K�я��|?�-�$#4��� ���j&��IHL�7R0������?<8t�T��V���m��$�Z�pD4>�rRo��h1Q8	e��O?�>];�q�\w9?=St�7����Ǫ��׺~��v�a�b*�6,�v��"[/��7V��G����D`�L/o�%}d��� 3C�f�4û+Tko�횏���	�M-�V1j���ߠ�ˁ��ǯ��iU�K�����{��0�J�����L����V���,P�$�0*;�(G�S��g:�J�KΚ'��4���%��8\�ם{֤-En4�5}Α<mn��N�4��o� C���vg�Ϩr�lfˣ�y�Ĺthg1�P$s����$�F'љ�o�T.#�%��Jt!��5Nf�EO�d�-�.��EN GY�� ���Lc �Lm�{�q��3a�Ԛ9��%}�Ȍ���S��M>nT��#%�&�ٙ�<#+��䜌!)y�np9g�6A`V����B�e�/�#�4/R�8���`��]>�;LQ�O{���:5��'�?�2���֦V�����*F(���O�9�^U������X�[��ݗd��v=4��Ŏ���}�OfK�ص��r+$B�*-�����J���p��:����$��,�I�����&�� *)���EDl���rɎ�ف�4��� �O��>�@ۣ��R@0����0�⧑ט���O��G��W���إs�"v�IC"e�q=�3O$2�`CN�O��|t�����)�UL:ڐ�!��X��b}n��a�l��g�����5�U�� ɱ�٭�]3tfmW�N�f�h��&j�-�A,6AiS7� 73�_�f��i4�X�CV�E���� J�w�r� ʖx+}�Y䂱����)��t}������GfG6�=��oAM��h���N�c�&t�2�@l*��׈�0�qU�����F�j��sA96�N�mu8N!�D�\�ޑSJ�;P�v=z߭.
���mP�r[*W,kbK�B�B���)�ú�7[���k���*���H���=���#��~�/�Ma.1�QA=�����=y_\��-�,ʺ	C�����*��|��hN�Gq�S�tr(8Q�\�;��g�u��3$خG��׍!�TuI`
 ,cx|��k �T�G�M�8ы��*�f�����K-����'H�՜��������n;���A患 ��!)w�Z�������Ʈ�moQ��i�&�q-	���}.X:��ŞG7$�����BKRc�O(�c���V��>��
���R|AK,�HbHc���z6:�I�i	�U@�[���2��E_��e��ʥn�@�>�7���zʚ.�;�3�{k�9<@�u���f����*xVv?Ng���߾:m3 ��׼Q�i.M)@A�~)�8{�/ �����v2���hε����h����$�ܚ���T���ٿT�}$bp��I���?�}���u`�d$�f��:�U�ݶ$ǈ�̐Xk.��L~���IOy�/������^ɖga��p(�6U�a�)�d��h�@�cav"N1��ý�o_Ѝc�p�rDh��K��i��sh��{c��9��d2h��ئ�� g;N�
s��3=��g�� |?��d(�>��u�����[M�m�)��T�a��|^-�v⥬��[U��LE��lz<0����u�0�@ጙ|�FQ��m
Z�䨹�>�E��KME�,�c�[/)ܘ���8���/�/�	�ǌ~7@����u��)���4��|��8+����ؓ����v��=�(����n�# �1
ߞ�)��A��x��|��ƏSrf������"hA)wp�8�K�n�G;�S|=��S�@Gj5��i�6����;����j����akEK?"��A8\��ʩ�N;�:�ҝ��dʟ����L�Q�����"�Wgh4���(����C��� �8���U�`îl�%��r ����꽋��"e�|Ot��i�~�^Q�ć�k��$׀N�<IB��QЗS���o��4_H6���6�ELd�f��`H��sչ�Ud�b��i�S�(5�\��Z%�R5�nܦ�I0CdY�P��p���ٙ���ld�;:��[yˮ��5�-�wJ� ������wL��+gŹI%���Ȏ�u��8�ɒ���x_t�C�Aw�n���_HT^��a,F�B��"ΙxTbvM�up)�_���0/����I1sǝ��4�1r�~B%L����U�
� N�-?�"+�	��%oM��g�3�P袖�H�;o7C7�l��Ϳ=�1�d�D��g��R�h�ýW@��.�Ѡ�qP�0�Y�ߦ�3��\�z4P/OC�Qa��W=���@#͉	�`����{����|RG`c@�M����^�ʌ>��b2�:�f{u��a@��@��L�d��=[��WC���l�k�M�SzW-�������-���5��?�VV����|%~�m]R�8�:6�#��E�G����&�Xz�mx'!�6k�qm�zc�1"�c����kc�A˻(}�SU%�3�˯7�w�KY�>OŰ�u`��Ac�ٚ)�l��A|���e�7��(P1��qmX��Ư �UE���?�ÖEy��D_.��/��<���H=w�$IjU\�>9nL�!� N���y�j_E}�xc.��׌�+��1�j�V��:����q�Wjp|�{<j_R��oyUt	/[��>�C�ںY@c�k՛�Mh�:X�]��-�[��R�K��T���G^X�8�w��Y��%*I�mC�+GPXEG^+n��y>4���v'�7s;�-"
�_�5�Qw�jʝ�y���=�����bX6�`��jCh�E��l��I�9��>$�/*u��E����C�ZQ�zko�J�y��eb�8h"�;��8���컠�/(�7��[�.�����8qV�-��AD\-�MX旿2�Kͼ��x	 ��'S�(l���)�@�6�C�����v�.�i�1`�Y^���D��(�1LZ��'+��Y��qJ u�<�mx�fwy~���A�Uٚ	����Z.Cwo�Y�/�{�� ܁�����0j�ȓԮ��1��:���:��m9\z�2��,>k�y�w�����%W����3����j���?��>:|�&v�e�R.��~Z��eef�����6WP$����|�	�([��Vh���/���N�~$���)�X���t��C��F`�8G�HQ��}���|�4��dE��O��r���"�"m���yf��S���I��+��ً�.|�PV�'p��"���u��I�H_�,������r�:��`�V�4޴�� �18<[n�)�ⳗgz�s�ٜ�i�oG�9�U�����%��s���n���AyPY
n��h�Ȍp�)��0�#��.���?\��T���1l��/3lQ}_�jy�_�Ƴ����c�	��,���#6y&�/�ق��&���gT#��e�*A�ф�#��*S�$��~�ڱ����	��8�?��&Z<�9��]6�N�Y#�HF�֔5tʰi���$G�[rt�k���O'{��u�ެ��������%�£�Vq�w{6���(Nj�b���m��A$��b��F���P��t}�^�Ж���5�F��'�Kf��q(rקv�Wۜ � ��m?̟9������������D�Y����Y*�(cL�j��0�G|tfsYy�{�TFQ��nW�S*���ZО*��Fw�����F�۠��Gf���[:$+7����B���������1SD��j9��n����И�Sla��/���B�mӾw`��)Y�����+2Z$���8`�֪�i�����%�FW<�L�%�InMR+>����ح�� SS{!�&���o�d�$��NGa��#�J���������|cC��-{V?��CaWÕף9zg�nxX���l̾�I.X`E���s����R�j���u�h �AC����5��m�'����	�o`��w���52!�ow���?��>}Y��J���HֽЀ��/�bU)�o7��ܹ2L�1 C��DP�>IOZ6Y���<�?yZD2�iD5�a��tṣ:
�F�?���V��xR���+�1���pHމ&_}�[�be�]�ZQ��-����qQ��j�Z�����3s )����.�5 �M*��4�_�x����e��*��!ʧ0<xOM~.�����ScMbUw��B���:����qL�^��\4��ۊrEʊ��-=�k_vF�\�N۟�q��Ɖ��P�\���@/|ՙ�c�����{��bJ���������+���+�Xk�w�y���̩&^3������"���V�`��3�grE(�`Ш�H8�f�rX[�Ϲ>z	q�C�F�_Ͽ�Ew���0�?Y��w�
!�A@�U,��u� �"R~��bFN�q�EɄ���B>S-���0�a0	%;�<(rh���g37c�	߰̒�*�LJl+`,�Ӌ�[�0�ٴLs�ྰܩ�A��q��M��AI��:��xc�=G���$ ��� 0C�1��D��+��H"��Pb�J{��H���\���\ZУ7W���̰"�t����x��j7�y�^)���ـ��T�'�͎�����5�C�$!�Ɖ�Ȉc���8�C]�oD�v,������{f���Ƶй�.:9t1p���^ĵ{���(�Oۑ��r�sv=ͫ���
߳�������I�p�t�u@[���j�;���"�\G���ȍ�"�%9;��F���+�b����]	R��ǌ~.=��
��u3�,=YT��hT���*u5�߽h�V��U��t��MlL������=�h��<Wf�͌�S"u��]�~��o�}���Ė�H�fM��;;�Gt=��VƐ�8W�'5����rS���q碵,t�5������n�δĐ��<�:�{�{��-3z���y~�L;Bi"���|N��fnv�R���2���2���5k��ȿJ��ȼ3і�ʅ˓�6�Ѿ�l j��4C���bb:t	P��(��?��`H���V]�����.W%�.���i����3�1AB"��:���:F�,�w��L�~ $ģ�qp��Y;|��
)b�{�6�� V^��=D��0�AJF�iP2���A8�
3�@�Z1`G��Cᔫ��(��>����Ŀ�P��1QjޙV�&�@j��n���dyM&�Q6��W�/�Jt���PW_"sD���v����V��v��G�;���t���Yl� ��S�v�#,�%��ң=��a	Je���G{���/5f���KLH�Tl1#2<f�p�����n���bUF��^X�g�����������8!�f�����a^?I��drmB�SX΅w����3�b��I��	8#�6��(-g���E��k�E~��C,���\	W�J�L"?ԕ����)����;��+�i�/dz!�mj'r�cYI� �\�a����%�v��o�2G����"'IM=]�w.�Om�#l%R�6b���� �2�UҌ�	�
X�fU�5(ғ7��m�J0y��.Eh��.�sc�q�N�S$��-���*˩�T�i!� ߠn���k}T��+�#�l&�/0��Q�@�����K
[���Y�f`٨�m�[U˘l��e^f���2�ݳ
�&����"]V,r*@��a䂰:�>�,�K�y&8�~�Ъ�8n�*n#�������N����Ff��SH��d���F�cL�t���
Q��4[ݽ3�g6j�)u$�7�#0�hu�ֿ��S�A�9�Z�<��C��:��nLo�B�0�6K���J�?`I�p�'�y?YV>\9/�9��j��O��2]@'����c�w+�mF�z�ix܏���eV�&�H���6��^劥�@�f�I-�P���|<#l��臿*�}-o%��ٕI�)�o#S�k�� iml�X.]j���5c~�S���b����^;���O&�xn�� ����u��UK�����(?�Q��
R�`�J:K�Ma�l��}ڤ��~��GZ�,�Zw�k4M���S��Տ���U"��3I�^.�9�V7Tx�ud�Jg�YROQ`k�w;]Ÿ.}v�y�!�QR�uC샱��~�)i��|�zS �7j�@���hi��,k9P��L��G� Ϡ:����_Np�&7��a�!�@}H��`!�� ��]��*ܒ7�fgďi�8���l'L�k(�
���݈�@r��6�T~����m%E���t��m�x�f�I�� �Џ#S~1�7�_бcQg�̏���v��N��Nء�������9�s�`-��80�?V�w��C�$����2EZ���NN�]�e�'�5�
f=%���b����\w��ϛLp*|�mB"��5!8��L��H�:Sט���X�:i|U�_ �M�D�-�gR����ki�"iu�Z����m�'d��:'�7�`z��SGEۿ+|�%���z���y`x���4��BM�V�q��@Ё�;v66s5W�g�ǑQ둁6 D��&��Ԗ�(��@4�N�a���U�7�L�Hs?�P�Z�RA����_RMH\7�VCM�*�ze-K��N�f2�`�fճ�6�o\c��w�;ڵ�0��+;���8���B��Z\=e�bl��$
��G˙��=�J0��8Vc#I�(����<pe
�
��=��E�U�X�J�r�r�v�SBj�n�\X���*�<�^���c��(�k)L=������eD��=bc�1U���E���g�����H�O5�7R���p�-fĈ�V�� ڙK}�Y��u��A�ް���)�=>�ӺR�����U�T���͠�ubj*���e���ŉF�#�_�T�W	��ХT�cU���Uu�������O��
�fۮI�RT�螅l�7�؊�JOW	0���zw���T���IrH[q��U g7TqW\4����D��1vXy�8�#����&�ݔ��� �%��V��I�ein-kT#�q�F"��~KtHVlޮ.����̇>2����*ʰ�;�Lԕ�,9��|����շ�9qՏf%o���Ddc$1VÛ�I�82�j��,	���d>�*���a��u��[��������e|�9�J�S� ��������	V39�,��;��3�n��uӀ��U�h���ٚ 6V/m�������!���V�mH���o��؝S��A�!�+*Z9-�爧����}"�����n�J4��:8N}\3N���ԷU~����mR�e��<�~s�ӭ�?ˌ�S��1P"�[M'M7x�R�^����VF��TG��n�C�E��݌���-�y�X��_^�/,�~g�
�n:�Ёl(b����o���n�RS����)�v��b�$]U;gOT�����ŢO�Lc^1~Q�ؠ.�[�C�UK; �����[oic�,��INx!�Ƀ�ɾUc��ȇ8�b4��eоȄ�-n���+�{��|��4������X��j/'9��41�9�����Z#G�~�P�eV���lz�x}c,��ﷰ��b���
�㛁(.��a��+|�ܪa7�Zo�~��<Q��%�Y�İ(���3��#���`�%&^xfƉ�1�)2�����Z��#G�t�0b��@�|���W��|��鬕�3JN������H�q8�dp��0F,��	��E3��UQW��ox��~a՘�l�t�{
	)����d�z'!�w*4s��鈄��(.�y�U ���@�2/���c������I�h��5k�b�ڢ�GX��>θ��9��Odb��l�*�R����Ku�ˬ��R���K�#Z;�Ix|z�I�N�4H_��V�z2��S�G(�uiձ�����I�K��0,�)a �fBRi����DM��_�K3����	���������ek�Cs݇8���o!=ꃘr�\��o����#oEc�3��^��h*��*E�l=5��8�WK���S�*����?�������ya&h��a ��\����Y��]�7wzt�BN��ѥ�t�����]��i��SGQX�<�f������j�������$,�:�xވb��P7A:�W$���~�����SUM��f�Sjbɤ�K�\�~��R�&\.ts�k���Kj�k��=�u����ҪJ�$ل�vuG�5���G i7��^�=�-�R7N� uK��^$P��W�Z�#��yg�r���!�� �ʚ��"��h��`n�W��R�!-�`tI�'�:+k6Z�(�^��l_�-�9�������Ȧ�.:J���?q۫��}��7\k���?9���p�8J��9��Ώ�ֳ>B��fu��\]�R�ϭ�����܋�AO�&sT�q����;�23x�ax�F�-��~tn�o릃=��Xn}���ٮj��p��|��w��kW�5e	9ݛ�U\c���o�|2".�D�O�ZR5`u�xz0�"�o=((��6�c����'N��L�߳��Kɖf�q�1�[�����+����P���1j8��s)Hځ��ִ �wS�������E�$�k��3=�}ʜ�4���~�� ob��ޚQP��]f�i2��j��ZTw8z^��G��W^�sDG�7�"hz������o��á;Y��љ/�T��z�ŮԴ9
��k���q/���B�`H��df�6J��Od�E9�-�m93�0�����Lnr�׃g���X{�" �hoH,���W��7
3F0JN����t�G�YT�"ڽ֮I<*��>�"�]��t�ΫF@YO�)��D�I1�V�=T�ϥT���?k�:��g��Q�t�����3=�*�җx����� 6�7b�cϘ�D?F��}�M�r"��k�}�!er�;�����Ͱ�+#-�w�K���D<��/�ż�O�����ָ.4�TX{��_�/��7k1���s�%��4�I�rw���괍��GK��v��r�Vsf6�B@I �#3��~2����NKp_-�Vq�����n
�"}� ��e��8[��kI�;p�5A����;^��u�v�g�0Xr
����%�40U�j��	fT?��b�q���^��)h����ctw�My��2%TH������}w ����%���0��D��E����f��?|]�^	�3��t����������~_U�v�d>��������L� ��>���ן_�\��S���ev��o�(;wK8��u�P��8QH���#��:Va%����� �A�~vGBt�´��������0�g%��GRob�IzV�g�
��e *��3�A�?�;�R��3ہqj����9CY(�[�I5 �6}�+�I	�S؀
���{�Sx��쎒Z�G��<��c�ve	s	��g�i�����i;�wjAw�]�����q�x~]1���+^b�^Wf����E
d��S�!�����6jO���:�L'Ľ�����~����%��#3���TVt��mp�Cz������I��E���o6��QHqP��eR��ф�{�w#xv^�D��߰��K�6ŦlK�F�-����SH���h����u�vQ�I%~:�e�vL{�~R���|K��럈M���lj�{sQ`���bM�٨�;Ca爾��+0{����C�ѝ	.ۼ�;���b�e����wAq~���sA�C�)�����3�jP�@L/�_+����1�Ty�K�[B^/ΐzgcg��aC�{���z��!L堬H�Mh�k9\{v�Zc9u�w.�S�@�;/�� r��<���1��D��nZ𭫁��.�^��$/Ӿ���9�DF����a{<2]{/u �N����{�5�Ə/��Y�k~* ��� 
���\����Y�e3�Ђ����A+ż�j��0�D)��`���4����yBZ<��{QgZ4$��~y	�\���ҡ���7��Q�G)m둥�z��ގ�`��?��h�^���r"�tP/�#Ɯ"|�w���g��OK�lq/��aiH��z��K�~���� ��k�xt�����[�(Oy�Vˍ�F�9��Z����D �E�a�x1yÍ�Z�ʄ�Á���2B�pf�s_�N1@�F�1���
�?�m�6;�6Ӫ�\�
)�j���܅j��͈z��h�p�\?N<���}/:A[
~� jcї�P���m�鲫���`v3���5����-@��0�܃���ͫ@�-g����.o�8W���R��V��!�/�⢧��)@}�kY�ֳ��[�N15��O$Nzv�j�,T�������V�w�[���-$Lp �a�8�#�V����*T2*?"��c D�b�U� ��{��K��`���HxB��=V�!_ȸʦ��u:;���7pAhk�i�s������I�)?,��3@���NW)��Ml	��5�����k�����N�X�'��b=[�� �yQ�Ծ2�qA�|��!m:KA"'�g�9?j�1�*�JW��Rq>�d�1��_Ҟ�>μ<j��@���L¿��vS*� jen�%�'��@���,z��E6���J�7����d8c��&����j�5Nν�n@:s����QQ�7k��0Yc�9��>�/*#�����@Q"� ����=�J���2�:(�8@��DZK���px���T���кL�QO(6�*w'M/D/k
c1ɸ\C��ˢj�71�vZM�w�����f�aQ[�������Ԏ���$ȁZ��1'���������0A�w�B�.W���sc%��������=�ͭ��z�XX�]%e�T����6������=-i���H)���q���v�4!���	�1�����ݒCa):���;�y��٫"��'�!��V�͑~<�Т��:2��(���r�@�Wn�F&����{\?4[^��6 G��ʣL�����۲�d����X�p�uNM:�.w�H9�+!�w��[p/���+/\Ԗ*8Q�w\�Z�y��T��zn�F��Z�u����|*�(|s��N7��J$�J����P�ԝY��m�[�hz�7l`��%6,h��PH����F��}cb�G�Q�Wq�Z��l��#̡?9�LC'�{o�aGac���坡�P-��Gf(��ǽ��^������
�_r�ej�"��7��H��Hӌ�e^���"��i48]��v��#ۙU�fS��7�;*@j����)��n%�?J����:ڱ�S�t�q��EX����B�+�v���&�̇��k���?|D�m&����i�sJ�eY�x֢_�����"���zB}�}�N<+߅�Tx�8$�4���oA��$���X�G����$�_���%f�D�@��6@^�ao��&����3ꦹ~-E&�������Y�E1
d>������&2�Z�\���L!�r�q�b��N��}���&�$ T�<y���������2?e{n��h4��oK~W�[W~�M�?�"MCu��D��A��_�9�I����\��JBo�C�f����0�E)
��L���4�&��K���N�]�����I/z�Hh�z!}��Zq�Y�c�j�i^���o�[��w��k�杯fx>�;��"Bk�2A� !ꧪ陆X�PN�d'x�N���Z���0�+�H��t�13�Nl�l�#��MX����^�	��|�g/v s˵�(� �6�o����(����#K=���"�U�x�T�2
$�YsС��5�j6_oQl���k9�nC1Ќ�\<�xe[s��c�~�MSH��qnXf_ips��Q�Alj��Y�����5u�5�I����)> �r�md��i�>܂Ѡ�.�q��]�P�h=SoR���ĥ�9/:
�G\�D��^����\%�=0ui�<������.Cm�?W�Ib9t������.������6R���
��'���g��²-Qw\`�v�Ɩ�h�����,��ɖ[µ���j��cQ���f.��+�i����C�z��l�hB���K-E��{�v(����2!��(��r`L�i1S�m����O�:j��[\	8іQ{�Е�5���R{�I��ho��l�1]C�7P؇S�Z�l����Y��h�4�����|��9�T �O؍}ʝ��֜7��rl(i��9ݶ�5��� (�a������p���/��kZVB��;���[o�d���>���/>�c�8K���u��p�׉	C��*���KX�bqy��)y����R%̫�PTT������]%v|��S��&�9�����FNzs�Om�I�9������Cʙ6B�d�f1%*�z��O1�b�R�c��V?����n����G��ni��]E�b�ykL��4m�1m�+�������J���]�mq��L�%��着f�Kk�1�[5 n�~�]������:���3���D݅�~�$�<�������=��O��W`+�i_#L����vP���ōD�ٷ+1]��e����[�I���dڙQ}7�D�\�ZH�wR���1
ޑ5= p� (�2�WԶ�^��XD�����?'�X�Ӽ2�o�f)��gn]^Pc�h�Y�O��k^��1DЁ]��6�5�*��̠��Gy��PU$+嚴�׼�tޫ@�&��Jn��������؇�D����J�q�Sy�"�L9b��ש賗���p�.Y�ޓAX�M�r�����VJ����!�Z�Ǵ�p���`'-<�M$0"���7m���Q��fݕ F��v�$�W�Wp����FW"�`�.7R�wn\n���LB)οH*�T���9��I(���{c�J*%�F�|�=>C%�D�����eQ��ޣ3��Q�cW��
)g����GnQ�8\؛�n�6Mv��:K��o?x���m���>��<�t�*�t��Kʬe�Eޗ��<
�q�������[�8ƾk�"XM�ye��yh�u!柤fc���槗Y[&���h�K(�kr��:`O̹����rcG x�z$O�IL��������qѨ|�'����ɼ�Q�W6���h��� K�{T��?�e��/Ho[/B���"���
�U"�>e�˔�1~�o�B�.];g�nb�8t!l�7��'��IE�mB�g���U�ե���sݮ��$��XR�h�t!��^)d�����&u��2d�$��9I�>�23Vg >e�"w7*>E��m���nZ��\�Z&Z��T�Tb"'�T��@҂���6�ɞ�>ؑ@�5`�&���5[42�1Qn¦�3\��1 ��:�n���Hb��x�J����r�qmt�1��~�"q�q��#ݱ���|U���VEp�֫���ka�����ζ�����~�AYs��Z�{U,9�d�z�~��=����:tOJ 欯�dYġD4P+M���ˮmM���/��p��-ѧ$���1�;G�g�fS�9�r'>)�����G�=0Bu�i�"�+��(�[B�q�0����kTՍ�ަ؅�=���O'o�RHj`��ûؠ��X��FZ�!Z�˳ :�3��@S�z[����B,�O8�����:>n�Ya^v��B]&r��N  ������VT���r�� �ø�UV�8p��ྮP?=�0�5���O�;��S|>
�9� N:�?���s�r�"��A=Pp߭���j ����L��Xv[�5bL�n���5:���,�"�5���-�x+M��<�d��.�ϯns�>��zUGC���+J)0Ӌ}��@~���yr���9�@�㶮�տ�,�RdTW���3���s��+��]!=�7�mJ�U��Q��_�m�\n?����\>/��6;�/j�X�D���7�x��G���bRY���Sʺ�x�#�L,EXz�vZZ�%������{J�VH�~�v�3[#K���Λ�K���w'�{
-�!�B@+�=N~F���.)���+=� �g?��@�j�D,j��s2M��^��b�-��hQ
v�u`���jz5�;���u­ �R+գ�ں�ƕ�{�'r���/A�l&-W�+K�xSd��e[�cwh �#�n��P��wۍT,R�ѩ!�ܢ�>��K�;b��{��'IL�D�,�'S��WB-��oԭe�Gg(\v+�����	���`�l��Ѱk���Bc�&����2�+�M�������������6��2�+�)��v�k�<�$��t�:w�����q��|���6���(b��ӑ�c�wo�*�t&z`��)Q#�k���ڐ��s����\���`�����G�%�;�qH�K�AȍIC��I���u,1M�X+��%V��0]�ggSKһ����t��u[�x����Bw)��`�=�y�6ǽ`� �!k�Au	1�B��()���_N'%�3�m|�l��h��>w5�^`��E�2��PB�P+�9�{`%]���߰�S��vV�t8��7�c��"�yW�m{Y�eE-�bj�f k��
�7f`�D8Xj<��������}e��(��W,0��"^O=]�a+��p�9N4�
�5|~�ML�� ��j������JR����#�,$��a�c�!��*���E�F�����+P��~�dHV�a��l�\����uܼ@&c���'���	��)������`ʺaO����q^���B�WA��_(Du匋ȸ�I��a7�J����zxY�
�N?�D��Q6K�'3�ڞ`�n;��n�:B���H���m����k���� ��3P2�˅��ψ}3G#'2K v>W@��P�jW�Q�\e��X�a�_�x��N�u]�����`8MI+p; ���XL�?[S�J���fb<��8Zj?1�Z�5L��5��w�=!��+u~7~�i�1��Y=Z<S빚���I�������;#��O[J�B��_����J������d�{�3�L�@���;�4�/�uX1ri��T8N�[��S$��+��߲Pl�Hye�[��cP�84���R�T+RDX��D<���դO{�o�rɥ��;�å2e�e[![[�(I\1,G��irTT��}���h��RMt5�Q��W�榆��Y�SCj����N,a^O��%Z��W�{�W;��J��%;�;�:�	h����)h�+f�ho�oV�VPwk��D�vc�K�{O��rNVr�ҝ�=H���B�J��&ᬊ'�'f5�3A7�b`<�J�X�ه/jM�m�A�����})�DVH��:ӵ1ڦ�AK"��0���I,�Y�y�����/9�x�+�,�56cI@�fF���S/%jG�]lN�aS�7u������ ��e�z?&yj! �SH�����a)��̀�i��kY�O�ё{�qBÎ���,�j�V#Μ%����;@�i#��ml�?�莝JO�V|�	I�?��.Zֳ�-�o?�E�7��)y$�����"�k�U��#C������ yq�"|D��oq��y0��;X�h*hG�b󼠤�x�.ل�>`��"�bZ�n�W�OU�sڊ�츃���CL�2G�R��6�%dFR�����~2���g��z�[p6(��YM��[�	�D1�9�0�
�!�=��ں��ln+ ��ao�y�0�Vf�5�w��D	����E|�	S@�����cc�.tD�u㳘�Pv�'Z�ɷ�	��'�&��(*"����V!�"��P��b>��3��))F��9_�6+���&�`��&`ݺ���@��wD��4�.��B����� �Cp<�P(R�	�H�����n-�-�*��-��؅�ʅ�P�.9��V���ݔ�$���e���K|�
�];C��cC*�����a��H���Q��Y�[����ʛI:
ꈍG�ן����P��5--ظ̈��B5�/�� YKAh�{u�5�V�o�_��������g�3Ɵ�Ã�I)�̇�2z�h�r[]��0]t�>
�8g�0<�_59�,���n�sX���H@��5�cJ��,�Z*Ŵ��%�i��<��t����!�fX�=ڭ;��9"4�Z{t
u�s#T�b��|�Yn+��Xt�r{�Q�O*��"Nd�2�g�;N���1w��<������#
H��L�d��aSV̰&�n-俑`��k��
��Na!��&���RP�B�-��4���N_�����6-'Oyd
�ز2����6�&à�mn�C�=��Y���v��M�b=�[���������P?�"�ȋċ�f/��jg�(+t$���\�e'֡��e����`N���n��۹.��t_~�cqI���	��4@J]�[����J�ڸ�XL(YY��=�1�:���Ώ-&Խ(R4���2f��w-�VY+�F�1�o띒.Q��%z�-:b��p���+y Q�|�P>���r!�_�@�v&��q���m_�n�f��%3�o[��i[+�o�ɶd/K�k�l9�K}��n58=�#��,7&�RŐ����4���Y������t�{�Q%	����Oz���$���'HՐ�䵖6G�ȆqS��#c��J��k�����B^��@��S��
z�j�D�{`���%4�:��O-�}/���;(�r� �<��H	�m]eo�-8�]dD���ָ[�.6=/eC�+S�����Y3�$�+����44k�'�h�`���d��� �(W>X�3 ��WwÑ�}��@��$ vJc�=4���Y6[|p;SzA`\��;!�;�	E��Qj��g��##г�ig��&�|e�c������Q�L�&�jҿEi�v
�� ��1Y0�p����ҥc�n�!r���$��H0�L\��]}Č�?�O�@aƤ�8��#�ٖ}%e���r^��(�,���6�ү���P���?�Z��2��Ŵ���y��"	�����n����ߛ��V*�"�Hc@��a��#�UʾL:Tj�����̸M�[e����C���0:=������΀V������)_����E��c�T�$��ڻ�����K����r!���ZqM��-�R*�oe���s3�����f���êi�'���_]e�tg���q6 �Õ�q�g���Q�<�������'�)�BߦZy�p���'�����V��f{:�~���E	e�gV�'���A�#ݳ>�8#V]ԓS=�d ]��M=x��Ǐ���Nk�E�C߈����������mU�vh�y�2^ɦ���f�	���w�ڣ)��n"��^�!�@���ı�������-JP��EX����:��{l�XY��@�=���KZ�=���W=�j"�G�?6@(k.�Zy���v�;����T���I��jꍝ��x�v8��W��5��ƺ��7�$�����oB��q����f�=](w��LM����7-�-�Pn_�����A� �~]�%c�����<��!r�W#�� JL�������0q�~�Ϯ�CE�r;���;���A���*�\<s1h��	��Rf�.���9v�P ���j9�ѽe��O����nIS!"7Kt�oq��`�A'x��*�z�4ph����7��'��� �=�q���>�%��c	�D~��쁮Uh���l)]����=�J�L�Az��o2�K ���6̞��i�n��E��Y�MpA���f��Z�z���˥1��_u��bCZ�]
m=�1'F�9��)�J���mG���(`;��p��E���l��9�K�I�c[2\������±��R�ih3�| ����m���@��YFߤ�ej��*{��D�8OV��}�~tqR�n���7cw+��C|�y6�xoMr�0/y����hs5����[oA{�J��`���0�ԃ_j��������D5�f���܅��^�T��gZ���ٖ�c���v������JK  ˙�c�G�0K�`���ޙ-=�j����x�f�r���@�Q����92ZD��`_X��YI��0��R���U��v_�wI{��`10��7���)�۬�{JB�i2�x�����ĩ@gj岫�u���_�~�
>�J��9h�nV��≇��>�A�l�YP��9zP�]A�͊�w�?v���NV!��^_��-�P�b;6x�`�S%D�z2)V�+�C��;���������O�x�BY�U+���YU��&!��ޖ(�<�q�Az�����2q�	o��S˨�vN��`�!%?�;~���s1����t��@|]�{�ZM�]�)m8��87x��fn2>��|8(�6�L��8 `��#�Ҡ��W�6����'�eow����Q$��=�E�ZL�_|p)0iAW'-$���͜�9�{+�a�������1;��r���m���c��|ú�����wY���`}p��o+�P�w w=�B��[�/@��+5a����ǳi��&w����q	���!�����Vf�X��)�Y5� ʓP�-�L_�QPB"��*y���q�q��~Ո~ťJ��_b���^��};5�!D�.�
�qm�������ǈ����rִK�\RL��${�α+�z1/[8.�0N=�C��&H��#&v�R�B��`QIFڨJE|���O��!��7����<mtbw�0r�|�۹??n����z��'H�^oh�q�Oc}Q�(��.^||��k���Ӗ�A-�g��d`��l��O9����+�H!ʾr_��C�6O���� �����/i���ȃx����y�Z��uw�d�W-�s�l2<�sƎ���Hb��RY*���y��[>@1��ϊ�^b����,�͞:X��P�BF2�le^n֪5Gq:W	5	1ȡ�JbMo4�5�coED��2%�~XEl�Rj���T�����A(��z8�K�@}W1H5^����W>�Y�Ϧ-HLJ�؟��Ұ[}jD߻�I�G�{ɷ��B��yfk�R�J�y��.���Zc��X�/{vV|Dj���:�����7��ed�NӁΒ��]j[i��T�0�8�"�w��>�a�Ԉ����z#�����b;̰�1��·Vtn^�RU6�gN�Ny�jP\і�~bq\h��5*`�Υ���Xi�����k$��A{凍���1m�)�T�h(/�\.ą�6��$�gS\�}c�=�zzK�b��r�Ky?�`2HH�l�}8�6E�����{JT�[��E�.t1�#6f��ݻ��T���IТ�Ik��8I����fL�A3+kT��L�'O<��r�W/�����������Z�hUrJݔ�|�J��:��;��I/OS�1�*��P��]�A���fb����KN��t'��lU�,�m����|"Ӏ��'�IRu��x�A�;����Ң������D��*R��&�Ȍ�s�I�9���IGdlX;�?3�a������?G���B���`��˫>�1�v�wj���^IBZ�l�Y@����7)�Kp�(�ho��I���)L�u{.��m'8��u�yhc��\L��lt���i���#��ﰚ�/D�/L�~f5��Wx����6���VP�kz���~�y●�_�BP��%M*nB(*P���:��0��Wb4��U@̿?H���E��F,�"�6��V���r��F�wm�3&�#�`�+�y�^�ٓ����wL��۰����/�gܥa� d���⨎���#��8�Ņ�D��c�"���+�y`pt�e�r4o]�wf�/����������_1?��P�mw�>�3�*޹��/ �0���)�RU��.�4��6�&lJj�6������p������;��F��{'6@]&AD�UHrcʾ̟�[�SM�^➥s!s���B����,�Xq��㣾���m�����ު���%�<>X	
���z	�`�_�b���� ��+rT���č(�Э��h'��	�ԘZ����Ì�c�O��nwIOb\_�3-��lk�P
[ъ8��M��C��u�ĴB��n�R�!��q�8dHn�9.)�!�'��`�#F�R�?��w���lp:{[�%�;��j<��W��X#�
��O1��<i��߫f��E̲���c�J��oe�-�K5VQ�H΃�O�Uf�O�y	��˿Z��5߲���Y��N5�i+���m��8��%m��͛�%�E��'�����{�H"6ajRa*]�>Pg�v-Ѓ?v���|�͢*��9V}z!b:��n�K�Ψv4<.�Y��.�� eS��U�^�vI�*R	rE�C��~9Ff��<(���Ishv�wp�2����/�ި��a���I�Yu]�¡���	>�2� u�M�J�,	4MC���ᠬDC�cc���Q����4$:s�%70����Ro<�������AS�Ě��˽犐��#���5�A����b�cyV#I�ҷ�s2I��o3H/(�W1p�d"��F
�Z@V���µ���_�1�\5�o����=b{�v�G��ST���~���lm��� �`�C���|���l���A��>|�o������W�>�ĻU��z
't�ڥ�;-+<�Hڔ���[�%�'@����]��y-g��~�,�H�k����:d��FW��u��Fg�|9V�����/�r��?%�RN��s�^A���BYo�MDJ�i��!�Ӥ+B^,�1Z�g����6G]��16>���W �f��j�aC1]W��.S�N�#顪�{���̡8ՊH�[�B��x�D��W���"	�ZhM ���|��&��W9d���=�$͍4�f]����%sc'�
�z��e�D�tl�V�p- ���"c�j�I��iDN�`�ͫþ}b2��U6[>x�f歹u�[R�'�`�o���K���m����aC9�78b#�u���N����T�rժ}��m|�nE����D
���D���3��{{0Bͳ!�)os�r�j�yw�	��C����q�]@��B�}��|c.�c/d���0�T@9�\�s�=�G&����|Qu�����`;c۠���
!3>�1�!�m��p�n�˛O.j_�a{��w&�`�� hҫ��n�a�
J��1�K�7`�!�E�B��4čH����q*�ɆN�6N�ٻ���ْ�r�6,�}����\Ӗ�b�\�x���JU$c���D����wm��L�,����yH
l���6�`�Y�Wq���)л��dg���T��Y[�;J�(i	��D5?�e�G/i�>F,��@<�	�/���fG���cjl�[����D�����I~��r~�ؼ��$/���讀�k+��[�"}�+�n��pǧ�����Rw��!�L?��/�imt�*q�W���Z����7�Q~7'�o���=N-t6�7�r��z�d�j�g���#c.�f���p��^�ti׺�ҷ��@R�C�����4�E�TT���4�0̼Vi�%�b�q��{l�\ªZ	��l�(�dƀT-��}�F��+73.�*(Ѩ���i��)�o�쮩�%�O������L��eӿ/��N?z]Lv�
��++/^��B��s�X�y���h����"�x^r�[LP�[d�o�0/xq��ڕE6��Y"f�ܹ�9�]кh�fV�#��Ŝ&RMq�q�\cVOǀ�8
���W�W��7�1�t����(T$P]�ج��S��].0�3�rǋD0��+_�~�OjorCz�!�	�V��)�Ǵ~���1r/�Q��Nh��Z���Р�-Ƴ���K�Pi�*t�ߏ���mt������5�m2k;��V!��w���a���у?ɇ܈,l/�75��ެ�wKk�뵽I��s"�N�(��ba�h�w5�h˒�F�|��*_Z{m�+̑u2!��>�$����/���-V��~ikx]aw�s9rE�X����ה����,q��+��%��DO���*��z�ə7���_#
�n������HO�<Fh6	��	��迨�O�?�Ք9��sx�i�8�}`��`�#����R�:�Z�����=b_H�i�O���
oP��2�r�脻�PL��76�����A��;���j_pJ���AZh<�,4��!Da�^sI��NЖ�p� �ÒC)�N��p>:t`z���-+	��b�U�l���J� �� J�Eny�Gbm+�=ȟ�޻��@��2�s�����<Rd�+��o+&�hƻ��
�9�"�|��}|h�gfPdVF������J�qq��/|���)�Q!�h}�ԿQd�$����y�Hx�a�Z�im�}R����Yscf�����1�̍k�v�E�5�aG%���R-��B^%��:Ȧ �	"��MJ>^��M
�{��:w�a#N��õ�ˏ٢?2F�+�%��R�	V�k�z�7.��SBQ��yR2�ԇ2�It������o��7����\���fৄ�JE~���2#�>hq!�mH���2��kӣ�JCG�슟�F��A�bQ�re�օJm$��Z�Խw*5�QE���[X��y��QLr:������A
!ԜS�|?��!\F�aa0z��{Y���E�m-��z
ſ�)�$ny���_Rg�xn��:��,i�O�G��:�_�@�3���:#X5��6���?��2�V��P7�
���٪A��u��6�LrJ�8}SL$L�b�;0>�?e@�&)��t��[�wQ�š��YFE桋w��Ltblb� ����5�'H������r�M=@����#�%tM���^1@���K�|�������^�[܌?o8
��
g��bC2��`�S͖�m�X��e8�{��@+��m|ej�����)�W-~L�-O�B�&��sL;n��F���yCu���ďzP��~ �W�l�`x�.�����	IGa��-�](
V ��k�%�V���f9~���Ƚ;Y��A�@5 ��Ѽ{TM�Y�C����ե4=iumV�UQ	�����4��ِ��
�q�����Jݢ���i5ڡ��]Wuo�Z�WD
��L��MY��~T�j>���5.�����R��Y���\��a8��G��$L"dz¢򪃌Xĕ�6���i�
hU��0����ԯZ�c��-ao�*q��Β(�U��u�lЋGˢ����̣f�� 9�E���:A̧fqV�&�8Xwo?��:d2L��}h��^lQgL.��ۊ0��|����0[4^�d��>&�PԘ�~'�e�W�u&�S	#��Sw���Y�?@j2���T�����'�|�B2I���Ԡ��A������y����&P4g��~���7�%��g#N9Ȗ�T�^qu�?�	�%ei�WY�wA��nS�{��}����$u��M8s���M����� ��8Rv�eUc4�A�i�3
�V{}�mW+ӭ
%��u��oJ��Y��9
O���,�x��YP����{5!�ּ`�]QWM�v���ԒI��m�j�F�� ΐ�r���zE�� ��:V��Ԃ���s��b�>i��y^SD�O�[�&H!�)5�/}�Ws$Qm8�Q�Rhs�b)�{���a�(9� ^w�#���'�+�9�Jt���ɵ��EW4��w����p.�{����>��!u=E�o�����i1J�^��';�$�����ź�r_4������H��UY=)-{࿰|Q(GA��
o����W'{�{$Z%Dƙ�i�����2�6=��f�ex��/ך�?�ټ5<�Ϥmffp[�I/�/%��mB�<58�qt�C߉�I<J�ڬ������ܶ�l�?J�0���L�VI�6-ry���g�6w��?��T`�s��i:}����o�ƴ>l�C�#:<��;�=�^�{`�7,�%N�9�3���pk�4�s�dJ4�Wf�^Yc?�&<0^0 ܁�I�g���򻏐ˊ%� ��$��.ĸ�*�6�^�|�6�5����m+gz�aȐ���K�p�MC�C������	���ؖ��}q����A��j�>����vޫ�>�c����Maq�Ds��Nv@ܾ����:�o�a�=J�|�D�� ���M
s �LX�uGm�L�&�^_��m�3C�J�зY�q�Mr�U��5՞�*\��Em�#���,����YG��1�Kg�@2c��E�r��A6\�x��t�!��癧�t��E��)���m���R�tд�.�W��%��S�xV߆��ر�
�>?�u�Bw������19ȴ�$8�߬Ⴐr,����!a=�����4���:.�v��^�܇��y��۸� �ۙ؇e͡f�_Hp����FS��"Z9C����J��`��ǕI�&^yF�y�?����d�ˉ����(�YS�f�#���m�������:��������!9�kX��x4�H��_�T��M<@絥s�֏Xq���z��
�O�����\F��k�L�5::q�$�$�0lY@��iˎxo�:�YӇ7��k�3�\��+�Њ*-Ϝ���IݐWR���c;��";�����@��شmy���[e�G%�������
�M3&H>��zv�5B\��#���Ƅ�/���D �s7�h7Kԗ�x�����#���K����ԡ%�X{ȑ�c���{04!OJ�L6���F���8l*6֛�6k-d�΀|Ҽ�l"��yˬ1M��:w���9����T" F
)�.�������KL��G�Ӎ�
��� ��C��V�pf(<r�%�Հ��SIE{V���ǲcj�J��,�G�3�����m�K�Z�ޖy��~(������_@��t�q]'5�B��=��Z�ۑ�?�|[<���i�O�O�,q�J���w��������X��VD`�֋+��	g�uJ������͕�T��,Ne��2��Ю�X�,��o�5���U"�>�y!G��*��!���x<���%��"�Q��^O|�~��|��(_��#@��\6p���� l����c����;��H��v�ݠ����y��/N���@^ď��)�;8K,~N�5r�	����Wuo��v>&A<g�Jն{�/��R�},5�a��]��0�5�S��P��$� +����{(�!G�I���t R�E��%���Ʈ�.�"���[�6ɴ�9��n�s�'�	�=x�
:BT�h�^�Y,����A�G)�.4�V&�r ��O�1�md�_�T�������Z2HP xXS������h�h�~}�]Atb2�}p��Dk�$[3*����r�^Q��[��=��K���}�\���"�8g�mk��0n�5�4��gQQ��z��Y�-Xݾ����M���zAQ(	1VV(��u�
�T�tgο���7��3�j�d��+�wEK&�{�:��u�t�a�r����!�!���.xv�XD���
�N����%F��>��'л1�-��N�|P$����W~i*�Cw�i?�5\������M���dU�� �D�����C8��q�)��?�L��R~=Ω�<�tY���#}e�*��v���v K��箛�e�F�y�dL��jdq����W�F
[��)�VT�Λ�$QnR���--�&���78fX��>�/}���L����iv����|�xn��Q\������2��W{�p�Le{wMߪX�X�:���Qk@}�!岘�N�r��hb�~E&đQr�J��0��Q�Y��}�ԣO��X��m �I��*��i��>�Y�:��;�axJe6Fx��J�|Qjl���S'�R$�g� ^I^��#����j��r��גAy�a���GU�^���g$Z�✀�K/�k���v�ב������I����vנV�?��U��L���2�9��]��	��L�;���Y#X�׿$�/�H}���g,�0�%���b�\϶P�G	�ˡv��dC:�Y�5g�_/k�A
��9���	9=�$��K8�1\����s�Q��	�x�q�U^Φ�d�&��WkrV�m��cM!8Y2�H!�;��z��]V?�j7�!�[�����Ow��i�	����e���1~b�ɲ@ù	x����^�7�0����lҋn�m�Y�*\)����u���ݰ_ӗ��p;��Mx��c�]3���9Y<'�:��!�F�`ŘI?hYr��� �'��TEN��3�1>�3�"�E^�S��X-f�S���t	%�,�& �O�y4T��f�p�~#�r.{�$�w��W�%���u�9���i�*,����,�L�J��8�Ш�rHA�I����xg��R�G�Э�e�D�8V����$�<���ؑ����_�8A�1׺~�]3�uV"��f}`��\�DO�����#�FEM����c؀h�u�8^fq=�	�vq�=G�mD�~-�����V�u)z�: �"���4Cr�=|p��>Y�����/n��<����0�/]���p�Zrf�Ɨ.�}�@*R�����ePP�z&Շ�@�dۻOѝ!����tqπ4|񡷛��J��4��������eHH����eHN��й��ls���)�e��Q�}�[m�栎��[!�0.�f��R��F��&�=]���z���{]�
y%��Դ�S�d�iد6$'����Aï�{�M�]#@�G5�6��y�=��(7!��am�X���㌶��)Fv��[�S-�gb��J�Ӷ��\>�Z�M_/_XJ*����T���d<�P�t��P�"����:z�i/&��`�q����K�1�6��c!���Qs��s�'tp�>� J���n�M��-�ژ��f�[�Qf�Y�0H'�Q{��a�L},�7�b��e&�Z���MЀG���l�xt#(���F���'N,�L�
�Ϝ�����d����m5�k��� �P|�MҠ��qs@a�d��rmpx�������Un1����] �'�� aW�g���i,=Na� EDbAfQ�Ğ#]�4�j=���2��E�i��K�08(��U�H{�^t��P1S��n��l�7������ҡ_�%�WR%�/�H�ߺ=���cKO�s�ZU���~�zte��P�m#N�4ҷ���J�φ'���_&Y�p���dF<�k���ŝh�Ti-,�PS#���3f�8��T�2�:�֟�H�j�-� �4����UQ���8�7%�0[�����K�����K@�0㋵˟l���ޒ��e��r��O[����l��Y��E�D����o��aG��e�,�-���Dy�u����H8��O�*��'ݯ-��ٲ�1��������x�����7�5ƥ��h:3���է5�����7�b��]�,į[>�Cʿ䎰��S1�c��E�띂�n�W��7�ԽUM}!�q�*�ʿ�e}T5����oJ�f�MB���l`~�*_eA{�����hWCh���w�Wjͻgb����M��"����J��$@��橚!�r��~O�]O`aᬣ1m��>�e������������E�@�1�ic��G~"�sz䞉ܟ=K��������a-�(��&�E�����3o&O�Y���O�#Jcx}�jBY�`�qr�$�k@��T�s��7��x���H+D��������SZݤ���rI/Q�#��d�.p�q3A'�(������)d���ao$uR:�f!l���f�l$�����Z|��B/=�:� 2�i؆�9��S�|@Y��������,�`�Z>�xm�vN�����8��o@
��9��+`�b���y-Y�&�E�&������.�)ʂ,����X�iYP�^n��7�ڑ�̄P��&�����S�LC,�g��
��@�
1��y�ތ}�aE��k`�a]_�AS!�iVk�x�����+#�n���|����v$���Wt�dw����?�Dir@�D���ۭv�t��>C1�dWn(�&��C"��=���=ęMA�[�+�k#�H���%�9�N�֨2e��d��:T������8���kX�Զ#�nϩgO�����`�\{��$)e ���v(>J�S�� �8ҁ����@y�G� �E�dp�>��J������!������z�Q�:�Z�QP�������>UT�.?��t1��n �Kh���9%61�h#|n�EF�qD�7g>e�"��^��j������z��tA�:����2	���p�MZ#����t��c��F�ѭ%�	T�yY����03�-��Ҧ5@�P�U��^��º���㮱e@�p3�Q�t2��$�c�dJ�ܭ�1E��{u���+E~���![ ��D@�ף���)9A!ts�x�c˰�TV�4��7�W�b��c��Ml@�ȵ��#���S ��ׄOa�O�z��x(��l�^��x�� cu�R�IN�&��F���=oĔ�g����W�Yv����L�?O�H[���c�x��[��c<;v�F�'QS�~%��L�D�Ҵ,��~��3�N.�����C#D�檞S�s�.zc �$���OI��t��I�w<��U���(�#\n�H��J~� ��;o��us��ԃ&y�v�sE*L�ݳ!bՑ~f��?Um��t8U>A��)|o��mg{������s�K���8�G�O�����.Fra��rI� ��8��'�LՈѠ.f�Δ�g�4�"bÍv���o���1@��QjV�����K�^ ������IQ��V9����Ԫ��R�B��)]��Kޕ®?l~�pv�-nk�K��"�-
V�$lS�p��W�r>k�6�u�[�2�>k���_�{p��k��+t)�D�~�����=��J� ��!@j�j��0���&i1^�W�/��7e<��$3׶���F� 8���'�vy���9-;�cP���#����72R"�������\Q���ņ�U.�n�3���Sx�n~]h ��u�R}l}�)�����ck��J� ��A/o�B���j��Ii'��������W�w���GXP�_ǨxO�ʁ�:��E�E�R�PKCK�2�[O�o$@	�����2Fȝ4Yj��"m�r��aC;0�(W����G5�
�d�wWa靃7F�g��^��B��c0"�L}*���Z@�;�
Τ�����ۍ��z�%/RϠNNtt�-�N��=8��;7g�+Ȧ���J���{�{h:��/�59v��1��DwU��2_H�oچGH�sU�������B����س�=�i�Si�:!��֙�mA�Б-`���H-����H���H�Gv��S]�K���S���Z��B)a�V�̯��qp��Фf�,��uЉ�w3����E&'*:��_a=T	�]�o��g�s��ap�\�=���~7���ϼB��uh��+�K����_��5g�*-[U/;�ä������t+�Q�N:�m�nb���+N�!�����[xǼI�-Wr��wX4��"�����dM-����Qe��/W�I��o�w7�G.��OB]d0�����_�Պ]0��ӫ�v�Ϝ��?T��ظ��5�}�'0��� �S�ԛ�e@IH�cEs&�X�;����0�˾z-��odUjq<�n]�"�8/��Na�ǧ%o�G�n1V��$�Lh�9�����ma�+������Fq�&�bAVY�&��w��PA7۝�B�1��:���n/q��8}��.��4<��ZyN�[��A�f�����C�!8��7�s�o���]�'��?d@k���}ǯN���9#7)��iΘ2X�&ɱ�Q���9�"OՔ�լ2|훚cѣ]�[�W~,(��Q��%s	儨��%���xV�7V���8�]�G�h�yPE��6S�Y}:�{��]�W�1����.��e,+K�C
�+�G����<�uR�u!���q����W�~i83���uI�T���K{K��|��O��ʙ��!U�	�[�o�N��gKmJ�W����v��T\ZN����n��J��pJ��̡(��<t|��Kw#c$��
0�ir#̑�A�Us_���Y�H�J��4�D<�C)p����Ȏ�SP���ǌ�̌AP��J�݀/��aVߵ2�Pc9�/�@�h�WA�$_& x�S��4-��nk�R���.�u �[�y�U�m�V��������@z$���>6�D���@&���Q�,��K��PP�y{r�����4n�6f��b�@_����eHV��_9�@��'G��H�U�~�Og��R��9��`�<�t]��d���o�\Z�H<I��]�� ��W��o�3ͻ�c�g��iEL��i���{R(�E�Dg�Mr��Y���\��!�#�J���k5�4a�|�0RblQ{���[P i��}�#�kz�<$��ִwi��B����;�j	ղ-)
���h�A.�4J�N��9���d۔��q�kf�4<��h��Q��c6��ğ��k�ni���^����x~�-3fF�tK��t���_{��î��ʊW�(A���SP��F�lr_��k�bl�A��$L�s�`��e�v�x]J$k�'�x+��h5�1mlo��WX3�g���Ҡ���/Y��#H�V�T؅%�x�L׿R�I��W���j^�QN���;h=� cGE���>�+��1�
�`>���m��Wά�n�A��l.���y��G�T��4�7������~1�*�K��[�9�K��J�}��6E��QH�⩱��8��!��懰�[�tC�ڰǼ|���6E<��D�Ȯ0v3��}����!5ۍl�ɽ��*���C��hdo�W��eiQ� ������d�I-c�t�eʭ�bw���7�7���H�;<C^����pic���側WYԬA���H5�[Ԝ����5&��e�m��$��A�F`��T�WU�JX�u4��҂=��=O�L�}��%�ynzM�B�F���GV��[�3�F���.���f�u��8^�����;3��/F���U�h��Šq��i/�Mh3b���~E���i�$0\�R��C��Z07Z�H��1t���w����S,߰vιJ7�w�n��B�b�1�3c���t����!f�,=�Ò������k�nH˽k��<A���B>�.~h�p
��A	UJ2�B O[��'`����5�J`W&s�V��:�3oV̹*\�c#�o��3o_��6�%;N��ȉ(�4��!���>�3�d��|��PXC���_���SG]�4��R���PN�-�E�P�(�B�fLT�W�(ee���_
pU�s~ E�c=-D�Q���*�1�ۆt��6{!L��$m��+�&���C3�O� .i�����z�o�r����+ml�K6|U������Ʀ��ڨ�qRztC@+չ��Ɍh��wĀ))8A"��@��m\�0u�|G���K@�0�����Wc��	d]2�/��E%`�_z5�!,�:�t_�T|)����ʲ�5UB�+�����^�{߫�a?����_�c�]��Њ�� �a@e��Қt�\��}�X.
���+�%Z��|1D�H0�7̑�f��q��A����O���Ů+�*��[���l�����c�Ӹ8j���N�#�E��甹��`��J]5�9G����P�A�)� �P
Tm��k
<ρ�`g�XHT<��R�?�k�̈́�`ZJqzn-]Z]��ظM���r%����t���p�4K��� vT"��I=YՎ*�|ԝ	�W��g�>�݄��xoV��I�W��H.�}��qit�ONi'�5�V�Ѵ�Ic^�T����
8i��G����[���ܿ�����co�����-��S}0d�{�6J{˾�u-z`{qma*%�哏.���B��#\����,�
�=���p�����a�~���`�gN�s�B��US�Wĳ���-��P������9 U=�*��ʶ%>���W~p�_kj�셉�&�ǰ[��Uh"�[�����ܽ�E�	e�dg@��\���\T�z�-�Y�;6��2jù�r��p8,��î\�KUhS:�;�4����;�OxYU�4��0�^��~��ZtА�&��9"O�GY��rmRX��"��و�ȇ|;�j"ަAsk�.,C�Q?�Β��Y�:�[��l@�y������sO��J�[7R	��N�jȆ "^q!`������Q���������l)��EuoD���&Mӕٴ�ڍ���j�EyL`g5��5z��Z;\������D�Ŵ�w	g*�)���!@�cD���˯��Չ)b	to�H�R��i�t_#n`������X�;K\�p�k�E5��]X$��1D�6�.N������Jm�^{&�ū�I�/Z�Rc�9pKD��{Z���}�H��aA3t���C�x�j���7���I��,�<�|.z$
y#]6Y�h���"h5�3�_Ł� ʅ!@oM07D��I�:�b�F�?#��v��,\ڀu�u₃���U�0Ԫ3����M���R?�3I���2��t��N�Dt�PD��^ԭ��O�CF�x�k�Ӏ ��~���T�X�4�����G��|;o����u�}<̏?���B��6o��z��)�*^���U���q�C㱝@E{���(���p��1�)�Bҹ�y5��O�Zq�6��Y^�������rj�.����N��f�8]��s`�����2q�\���Y�Q�^���nA��d��pɧɤ*:��h�)�W�'�Ż�j�I�"b}�����3���[r���];׋�\d��w���0E>{\����3�e"�"h{f�f�2Kz�{v�t���JI���-b��+2�i\}�[���>��b���~�嶚�8G6�F�!�D��}��Q�yS��a�����]���S�5��eC�k�h���S^Ù�=�.��i��yL7.�C�$��E�/i����T��^�
鮀#o������G�rכѬŉЉJ�p�6��l��o��䶤Wxd�~� �֔듼V'͓_�\�_#��'����N��I67�����B���By2����~��){�v����Td�l�?�2J��	h�e{�	��9%��$=X1�ƞ�o��Zf��h��)M�i��.>�'�ࡎ3���ݟ��%+w��$�oi�#�o��5�E��f�!xw�� bVW��K)��?\�ð׍���=��m,�������8SXA����.����a����CP޼���5@U�%`�k��fI���wĦ1�R&�ua��7��𧵿�#`�"�N���I#�i-%��O��[㭑��)$�0�+vq*ODw(ڍ��|���tڝ�dz�j�C�٘"��	`L�I�kx�Ub�m���L}�o��M�ϝ�l��s���B;�6�7�(^GRJ;��v�Iށh+�9��r����,~�^�>���mRN���zX���IU BϦ@����b���[��G>�J9��g���B��	�$�{�y��=�2��L�H-�n�b肿�Y+�g�\K����o&k6(�.��0Wv6��n�уN
z�?�=��	���dQ���"�T.���}����p���D�0(���_mѤ,�Q|=f��wO��Y�|���� C j�O�EȾbz��g�l�B�� &����r�	�N�M�O�s���y=������(�Uؐd�rg����fm��]'�x@R�iG�V�о_�*%�C�1�S�M9H�?C]���%]ar�:lW�Q��W��$m�.�*y�ai�Gz�ۢed�J����ǍˢJ��"��d���s"-��$T�ۗr��xG���85B�C��Z<�f"�b{������ �Ba!�J��rx�@������\<*o$��=��÷h��+l�9E:��:j�L-V���_���w	փ�K�ۨ��'�f�5�$�tN��kx�J+��$������Gq��1|D]���/
�5�t�V�2�����Կ=8�VSmT�
��f� d/�+,�����rLq�q��x�	��V5��R���+�Y6L�5�Z	��G�J�K��(�3�|}�g#M��Gv��Ylb���ʋ;tݓh������2*r�9�n�(�.�,���Q-�LQ��2��u��&�Vg��&����n����3/��h����J4R�����y��4�:Jn�SE�C���үN��ߊ����H6n��+n�r�K'	�L��xbп��&�,�o���7�����2G�K+և���Y9����y����m.] C�@���t�BS�f&�B�P�=���(�p���!D �ރn�ɉ��_#����p�k��y<�;�M�eh�/i$��$�B?�>R����^lX�8��*Y�b��8+�oc#~
E���x?*gt�/���9���P�[Wb9��"�� �֨~���?��$������b��b7>������kZ?Y3zPۯɖ:��YtF�	{1��4�q�{]�D`�Md;,���!Ee*휻�S���-s�CcK{�M듈V��t������7��w��w�Z`���d?z4���`�qO�拳�n�͉���	�Qc� 0'P�2�\·�h�!����5�u�6v*`��o�+O�����é���H��wc�1]��n"�;��?[ɗu�m	�G@[b4=CO��`<ʣӅg	���~x���Z�ӽ�W�B�~P���-��,�c���݊��D��+a��2��	�<�p��A"9N�SW�c��S?
[�MSP��{Z7�^�\�	��ʓ�P�ʬ�/�M͛Tk_>�^nАS�@��S�GZL-��=�s�M�v�`:���q}��R�Ip�%﫢,&��V��n���n�r3�0������`ن�G����)���o�����j�<C��V�({MSc���7�7�H�a^���x����(?�i3�.�eL�p����h�1\?m�pd�����f->����#]�,}{�ט^&"Bc�gؤ"^&+rp5"�>Q%�ό�y��#;X�6���
R�<�[Z�F�Ft��u�� 'e��&0�/u�UgD���W{KA�k9F��9����!LR*�T��v�K/M��C�n��v�����qϪ��w�,��Mާ�E�>�)�\�ᬽ"u�f i�˻���W1�����@ɗU�e��Xl����r7��#���¡�#�=�(��_����K@�{��B�r�B6�����k����s-�(���yf����F�k�L8��[��k��i��Z+���N�	�&Wt?#�Hmz�6���O����	�d�Sb?��æ�N�LNRMw*I`8�8�V(*��]�{���+_*i��&�?b�z<K��I$�vJ�"y�nTQZ�G%� p�]
Ѱ��ޝ3j� �
��b�=�c��Ϟ�����e����[b<v7Ԩ�'�~��q1��ģ�?�*Qy�W��e�q|1�X�$����y��^	�3)��_�yGfǝ	���h\YW�gE:��W���g\�s<֞���G�by�7���C
�`����&�t%���0%��X�|��E�jP%�XWC�_����8'��w���7��rKϬe�p�@1�'vIj>w�A�z�Ddڣ�f��	gg&��5�����b�Ywk��￺�1��y����	Z1�*lz�t�Ʈ�S�eY��������}SnPe:/!#��^�v��e�J1Gv��7z��|3��=��D?���qM}|q΄��f��ilۺ�ZY�$��A��`^�Q5*(R��]/>�@Ҵ�w�v˼��pSz	���V�g�I`=�D��˓X@�QŸDz~V^=6,��8x�8+~��}"�%o��M~g��΂Q��\l�x��H����[i�#�Y���Jh���w��t�����p��4��)�W�L{hm}Z��]f��TV���b�NkNg�}-͊�����U�+v�)��ņJ��k�?jQ�#�!٪� XyBc���h�JC�I��� t��T�d��9�n�z�����$2��%~ �^��'�YOq$�şK�zi'��lvle�uI~�����q��z�>Aތ�,��I��V|Jň���tO���B��l��98?R
$H<q�T����>��Ƕ>�T��*݅`�r�㔤�Y�H����^���v�'IZ���$�����vtc���J�_�X��?ę�ea#/2�\k��?)@�������.����$�~����>*�C�Z�Z���Y߆k�g ��i�[�\�r�@�J��^���x�:���%kz!�+x��tg��碈J�Н$�5�C��9�1� �,�f�qt��7F �pC,Y 0���$�=�y}���1L�1��CP���j��b����Y	 C��oC�F@|9��[3�ȥ&�E'�0$Ț���ij�fJ�"��Y1�.3;�Ӭg1��m�T��e�F?lԥ�����)�;����R[�	^���Y)�@�׼������N#	C��q��֮B)�	R�h<��E���s�*���b���
	�<�4�CZ��1�G��U�"a!������m���c7��{`ÉW2�3�s�E�~�&�kOj��Mz��2�㗟��)I�[����-*:ܣ���m�|! b�pj���) �Vy.R�FҀۘb$%e����i��E�-�KD�zT*��ws��)X�u������	n�CC��E\ ����}��5I*;�`�#����::��4��v o
�YVh65�S:���6?.,�"-ʓo���8��!�2y+O䍴�T�0D����@�v��	�-�m����B�s�`���j�`��
��?���:��qLA�籨P�%���w�JBO��M�e�ܑ�3�fU�yV@�t��[�l��r#ŕ�m�g�vd'���9�x��]|+:/�-b沠�r�ì�R8q[���jk��cjGF��R����0�$d�3���ʗY�[�xN������3	����͇�	�n��Y�Z��H�BJ�����Ƕy�g�	XW���`<A��
v�.s�M�'���os���%s)K�x ���1ѱ���tr��e<�L�n�I����dȵ#����r>jC��,G}���U�+R��N����ݍ��&x`^�F{
����W�����X�QX&`�����:�t�>b�Ӌ�e�k�	�t�F�ܷ�]����H6����#}���ɭ�A�Ն\"%�A���(? eLe1�#+���vo�>h�g���og�����c>�ހ!��kb���OLY.yZ�TG�P~�����QNp�#����,��0ƴF׾a��J���6@N		I����=�5hK7��G@��W��.� ���I}��Rӫԅ�:PbjR�����1�p�S{��c��Y���9��z�����]��M�1M����0T���m���C?<1rW\��r��A���(�CW��� �.�H�d�+ں��9��F�`/B��h���a��LL�����t�Y�:͐�,x��z��>mFΗ���O29��O"Ea���r����n�������`?��|Z9N�jP��F��eR����`?d��EP�q�F&Q�A�X���$N"@y)�=qP����Ia�S{v辈Py�6��m+k% �@�6�.����e��oIM�������N�!��ua�UZ�4�}�G7��"-��b��K�`�T������%���+��~9DA|�PFZ=���}�3s�FA�UZߖ��A�eh���Q��1��*$�\���xW������ݖ���/��ٶ��Q��s}� �����G�����|0m!���k|+oMn�K�rP�x�&T��o��f$�є�����kn���b���Vf�#���,�!���wp��5F�_N��\�)(ά�
��2������$�9(��1P7#\�f:�\ÙF���%�w�(��앿+<��39/V�B'�=ܘJ\^���=�tȌ�le��d<VvT ˳�'����5��MF-��ڝр�|G�~��D��faQ\:�c��6�_je �5��ZM��Q[K�q��V
	��]�~���S��	E^&�M��q!ۅ����$4o��5UTm��e�in|�yM7
�d�a� ؐ�1�uc��\*e�c���\!���Z�%�|��dB$��HG�~'�H�M�`ZC�����Q�=U�G/���j�Ik?Uc�
~��0�e!�,�_���Һ73z�l&�6�c�]���?7q��=�hi���'��t�Jça�IߪP��*ݎK�.��� mT3(��F�w0	`�LC�`�x��Ҿ���1�m���z���:�o@y~1�&q�q���Eb�q�H_r��l\��
D�]�K#�VŽ�#���VW�խD��ОkT���9Ω�)��=4G���^����!�`��A�.�8��㵾+n�"�? F�7����x���"K帰i�t!I`޺�t�)Ƹ��� ���W
d�_,��Y[���Tzd�n��i�b#�+�2�&�1�a[~ev�0�5�%ㆹ��<C�T<!��1��~[Gm�K�xc%��!���[&}�yp8�����XHrV6���>O��,�!��4����H4*3��(����i��)�A�	�F\h1(x�[�C�
�n.c�US��f>8 �L�ޞ?˝AGȭ׬e�u����j��MQTM�J�p�>$�z������w=zm�C`�>�nJ�}&B(喘���Q'���f��9(sseUS3�(�3w��Wr��M��C�D�b��4Cr���>=B)��|�/���kmo���w��H¿������ 4r�bmUk�t����ɭ����rr\���6�J��ᒂNlzCu���e���F'J�i�a�r�A1E�6�W�K�EE`������/:��mߨ���h�~�]��9���8OA�mv�)���d(l%�"��Z�.��m����io�镧����{�ʣ�_�׮����cr%>P����5�q!o��4[㐺q5v_��]�vnb�b���T0]%7���*-
�J�=�v�Q�ʬ7��(�Q���I���ayCTg�I��	~?XL� nWW����υP�,�"�/��1��=(��@������4В�h��8�gph6-vq��VA�j�&h��}X��2�U�L��
�{��=	4,a+�u�%4VD{�l�3Q�%Tn�=�o\_���k�5�+U?Gt�m؂M4��$���D*k>uk���Q��6�e�,{9�M����q(7�V������ő���3���h�=��ڗ=�Ա�W��[<�W~Ӥ	|6��G�|6%����R��q8����3nt���d,��H�8���C�PЀ�<x�-�����̞B'@%�?28��,��j	�H�O�f�:�i�0�A�;'�����.�V�=d�SCgM��b�d��s)�"��`^��*D��Z��[�|ՎS�����3��sWK?���O�|}]@�/
�)��a4Uk��(Ѭ��"���w�X˕���sx9\��(I;����/���ڌh�g�?y��T�l�%���X�}u{���L���������W��j�Qm��7��`R0�	���Y���Y�U��~%�#e��)#5��t�{���#Kk��~g�?���q�|J+?
�-R+�ty"H6�Ʃ�ʻT�y����ȳ��e���ka�@�����������-�?�c��P7ќ厖�
L���[-��6e0s5v���w: &���KH�^����n�'��Ίf)v���f�C>R���L�����eQ'osP�<���-�B��S8T4 �ʊh�g����a6Ұ|�W�"(�w�{��e��}*x��e��_V�(��De���z�6���� �%�A�/� n[��<��H��֭���'%�d�9���N4ڊ � ��%�^G294x?�fȬ��
�D�429�U6��ޘ�
��?Ey��¸�):���՚��3��H�ŷ�N�)�;���5a���\�$d�Sy)��+�j����+��3�c��`K�L��c�*o��0� ����*�[Np�J��yάXt�=��jT��m_�y���×�m�P���P���{["��$�}f��#�>����}����}9n�6V����Ѳ��݈��j@W�̡6�r������r1���+ޏ{S��ٻ�y{%��v����g	�����&��I��`��N=�9
+�\���o�� ��[S����D��x�-8��z�nB.���&��G<c s�]��R%��w8�%2Ҙ��C�o��L�-X����Gs��r+\��HfL�����V4��Q:Җ�&൚�@���2;H�𽉖e��!��$���xB�I;�Jd���˽�;(5���[�pܠ�)a0��(����l��G�ߧ�����U��!,���#M�m��L�yP�C4��?�b�߭F����-Q�5P�]��H
<��"�yf~Jg����P}�]Y~b��q0�繗Ypc�C����0�m�kt�� G9�.�&���k,�H|��("�*�w�>��aPO��L�!P�a��^|�����h��ZiB�^�T?��C������ɢQ
2�W?,8y�i�����Ģ��h7�&)�!Mvc���i���|����|�T�v��u�X{��Q��������n~�]�ć]>sG�h�'�<��3���#��45�5T�����-㬾��� �d�;���R+���0���O��	w����P����5-X�$24e�(K��������U�U�����#�C&<��	;�s�xi62f/'���(V�zHk�\/	t�c��`Ҧ��ZA���2�qrQ{�D�k|�v'gn�tJ'�Lƈ��t ����0� ���Z?,I�4���W.鱳��V�a'jՔ%ͧI����Z��1˧��<G�}��C�[���
��H�sۤ�@���E]X�'{��|]u]w�A�S[ɔ�.}]ȵ����>���6�|�n/�~d�u�*�
�k�W���ynJٝ8_а?�Y� O�pG�lJ6���8��uzn7>\͌6$��[Y��xe#IC����gbO�m��ۯI���/_�b/zqc�e��@���٫&kĿXG�4ꅔ�2�^FS��6j�E[�1�4
� �@�$� 2J�c����(�|ۢ�w!w��본4Jl�5��s� ?�;��ۇ���xh��}���p:�px�������E�ÿ��GO�&)60A賓3�c;?i�z�L�A�;�����3��H����� �q���0(u8��,���#G,�Û2R���s��ӌ��4�8n9<�#tuJ�v+���"'�'_r�(�2�&Ǭ�Ɛ�W�5s��d8ٝ�I���W��D�K���p1�e�KLR�}`j�V��PH0 �V �i�
�^�'�շ6�w�ꐾ�
!��5�>M�GE��.����`���~��ދ)���O���S��).�,i�!���t��9oamﵧ���8��T4�1ɗ��N����ū�c�Mh�[�M���S��+q%Y�����i��[��#��_���M98�.�N,\5v�����'���2����2uǐ5��(���P��+Z�'�;*M[#�%|�axx-�V�����KGF�B��G��·;V�x�}OH7mn,R�_��S k��7;��������gq�藴I�d{�C�/o��F�^8��~l�l�iJ��D^&��ݥ}��Brd��������L��8�"5Q�h�zD��,��� �������?>� ����<;�r��R��{�%~���y/�)��yfT��µ1�������3޵u�h��$���\�iw�G
�ˣi���.'�!h@,��Y�������.'E��^}#E83���ےX#]Yԧ��w,E)���<Zֱ;�Ѓ���� 9���^�)�8�z�?�(����X�w���g<�b�������w��>1���V��ZM|-���+�I�)a� e$�Ato����1��O�//�y�y�|mh(#����(��k��`�n�r�JJ� �#ƚJ>��S�L���?aٙ�2j�}��lnZ�v�M3֕
{qj����?U�Va�9��!�� U�BM�q��V7�Yy�p�Z�{�~�R<�zRXVfec̈���8G���o-���
�'�E}Z"QѲ�$�&�>���s��h*k�ivM�����k^Q�Ϥ�c��C�1�	��QY�v_<�)&�cn�Y�I���6�]2K3���MiN�F����\D���⠃��_U+�.��'/��s���#��_/��F�E�27u@���b���7lQ���壷�7l����Ծ��Ղ_`�΂�����!��b	�\ߴ1"�V �6�XXΙ��	�Z�Y%���F G_n|@��NZg���`����%���ٚ����ŵ�!�3� ��?T�u�aO"{a KQ�����@��@f�(�=%2�Z3�3�&j�@ θ�B3���^��	�5�J^���̨�������TtR�y��)+���{4�[���dS�)��ϼf7�����f�I?���4��<��-�G[�4�ߩ�Ǹ��p�s����*��fN�������CWǕ�=]8��x�+;(�������ZC%w���f�bbLPYc�9�ꪼ�b.���t��L�\��h����;m_Y5g�J9�̇���ba%���/Sؼ9=��,y>��/��̨�J��)����Ƿ���F5��r��֡�:�*9�iJ����΅��>D�P�o~���@������,ɪcO���M����Šy��Q�(����5o������P�(@n�� ��B��oC��vOp2Xz�t���?�琻�`���U\���Z:��N̝���H)�??� 6m��h��v�S'�	�a̟ �R�f�)����D��G�/-���q���)g����W"�a��F�4��ݵK�G�n^�ᇵ)b�[�C���e?і�"e��ͥ�EX-z?�y^j�j�)�T ���<�`.w�º�z�i�	�u�A]��lF���8 A�F8촣���]����¯����#�7fG���o�#�Up��ޜ�T<��y�؝��g>���gp\�J�����������&�&V7F2���TIc�-�CI_K����no�\�_�i�e�X�0����pH&H8�j�HLwc�p<F*p<�{�ˉ��M#f����|_&���~�+=�@�r7)���Ѓ���-����M���7o,�0f6"�|�E(CR�5����s���r�ľq��� ����sE�	�T,�� ���c'i�9f4�9r,���ں��:tL��VO���1��g�=-�܍����UA��娑xH�zI��P��-������c��c���}j�%-�6�9r<V����Ǳ��@�h��`*��V-�o�N�̥�#�Q�@S���:�=3\�[F�^�Mn�L�f��f��7++��h���pbA�:t���U��%pl@�#z��\h��tO���{L�g��94���s�q[y>�����p��b����h<�xs{\��ky�������9�x;�.�тs��eʓ�M�	ξ9��	l]�q��8[Ǡ�؞�g,�����{W�y�/�X|�/�ܧr�vc� "�3Mڕno/d�c�A�I�qV�E�4�e`�]�3#v z $���� E�ߧ���ϴ���ԪpJ�h����0�6�����F��	 ��墂��I+�Kv�K76�m�ߴ�ׁJ�V[k_2[g,VW~�YD!��}���_)S��h8SP��l/�H(���	
��Y�(� H���m�j�����Y����p^�*��)O(���u�'��U��z=���|�D��M�)�6o']�]��ܝH� ��=�W��Qh������g�\1�ͫ�u^-�K]��UH�SUtY~h����D�����f����ns�,�H�D�6~��v����*'1θ.��|����FXF�Kը�֚x��m�jh���^{��(��O��ge��Ʃ6^�`�T�UQ�JCW� :���Ea�����c�NQ�����^��I�I!V�umHR�뫡�QCf�*u�p^-� ����CG�託�3\�t	�^'����Rq����J�I��v���]h��d�uM��Ts��P����d���Y��Cq�����΍���c���Z� ^�R����	�
�$���~���]��e�9�{�tL*����.I�)O�����E�}��Ց�)�����	�Pomjg�7���t�d)�f�\�x��`��_G�o���없�s1�������{��l�s)ǒK������M��� �R1Ì�S��X��D�"뭻Uw������>J����R�R�q=��𽪱����ܘ;I�$�q�ʐd���!�{�$��xJ>�1�Y�/T���m����=�zg�<3��;�����/�b�a����@I!���{��q�>1.Hܤ@}9��R�vQ��,C���T���P�;��7�3am���]��6!\����ôURV��I����X��k��˪[��{�©�	�:[�5���G �H���-,l��N4�;�U�,�iM_�O�����L����&�+ֶ�,�[����҆0�����*K��n��$����)H$X#c�Ts�C�֓�� ���PF?����m�9B�ol����6-���6A�=Q��9ۘ����L�Y�׬r� 7-C}�δ����#a7� Z�@�8}2�k
�
<O5��.B�������0�L<^�͖ڗ��j;��E��#ѿ>�l!��H{����RT�࣐��e����WS�Q�y���s�T�����.�\����>���V�T�=����we�-���kQ��
���$|��Ce��{�^�,vf��=�N_L���}'U���L3�g+b��$5ש_�4IU[!#}*�3Q�k X���-���U���M�м4��Ku*lz��C<�&L�j�������rԞ/�j9�E�d���R���S@�[����W`җȤ[ە���'@*h�i*�HR��8= =������<�_�/�2�S��a���@K�n��gм�����Bd#��s�J*睰}K���m�3��*H&�ed��،�Yx?1�ɌVg4���I��2{�<_hŘ��i�h+f���%�[�C�9� mK��CS���8}מy�=��l�Wtt��E�(��f���-��l߃�61�j�WzD��d<�����=�\��#�
�(V��ch�lӞq4>�Qk'�^�ȳ�8�y6)�y:0*��7,�RS�;��6����%Px���|�=�g@ ҩr�T�FH�ԾآyϪ!��f���pg��E!����E�t�I;ʩD7�FZ�P{�8*KT͏��l���T;1�L�&�]����
�Y�\�F�+f�e�h���:�1K_�%������$��KA��,.��}ٖX��G�y@"���x���&�<����'�?�N_
g9n���Jb)#����[������&�.�7G�*��� ��)n�[o����Z��^�T��Ĝh���d����� lI����<�^��uW0}B�O��=�/ǹ�?/��8�����-g���NE}�R%����}H�ȵ��M��h�q��ѭ�4%��#%�ؚ%A.�4��]�/�	�Z�i�K;z8$d��6���t�*��a}���7Nށ��k�q�'�Ks>^(��fū�Db�����S3G6ꁳO%���y��;"�����(��|�d�:��rw�e%�L�����4�Лt5K�k9/�E��]�i1t�ˢ�(��#`����k�"T_VcgAB!7�B����g(��L�;�ܢ����h�b8�5����TC�$�h�x/�����N�^���D�>�՝}̒�ˆ��v���,|��S3��O�5������*5�Q!-�x�����Ő4�`�0·�j+���ƃё���%*�旀��L�0�BP$B�
}�_�Q�����#(����ɜ�� 	�ܒ��MI{1e�*c�+!�Eb`;����*�ݻ�8ѿ�6��F�*>�K�[������ 3L�^�n�$�pV���%�Ov��Ill����5��Gy�b�C�P���uT�1��K�Qg����B���lw��d���$F��$X�[jV�	�#�Ќ��Y��Ë�<h"?8�2׿~m��M����WP:�Vyg���d�p�/�Fa�p����tl�Q*˝�Z
�*5���S��O����T�]۴�X�
��+fRc5}��_��ĥ�7V��)��+PDЭ����tՈ�vG*��kD|��%�s���v���b��G>(;귺z�3S𪬝���7bQ�\���wdV�N\1u�$Ph�̘�h�v�:g���uT��0���
���!�U���^�y��=�ۙ8^���.�sQ*%����)��q����Z�ֶ C��dNvW+p�*�JE��R��wU�܉$Z�59uu&Ý��.�@>���cAl��.��_�n�G{�W)f�%����+�@`���%!f)3����~{�~S��Z��5M	C����kF}M6��-��06�^�1֥�(g����T1��}�2�ʺz���Y�(����hW�0��/�P1��n�N �K�iN��N��GW���3A4	qg�A?�!���eT-R����<e�R9^��hXem!<��1�ϐ/qMav�+ņ��^=��60�"4Rs�jŃ6�r�Mǯ���Sc6.�2��5���b�! pA�X��"�.��%��gB9��@�Q���θmi.
����@��G���YMh�	T��4��?L�~�0��~f50����MɊ�	�Ҕl�0�Uh	�9��-�o��oQ};���Q�����������y�_��+�pY誸��T.�������*�8��x�3�o�%���~�YS1 �~qo�U7+�xd�E�ˏF�T�qy[(���mA�]�����_��"�]F�u�	��	�5�PY������2y��52��t�ͳU�<��d�Gx�y�-�c�h]�&�H\�d�R�<�ͅ�r�=j�)�ǰ��X�\{����aݍ�@�l��������ӂ�0&��L��Jr:�{�~�@rÅ�h��!�P�G�	
�,ۯ�	Ҏ�k�uE�b��iǋ+t����h,N���Jի���to)������ �b�����2�,�W3��\�ª`7Y�߅tT��i�׊����mնFoRD�GW�G�l�:�ӿo��7��x�&Tp}�p�ٲ�Ƈ��@}�i=��h:�ߌ�>,�/χbg��XU� Bs������V����4Q��E$C��[A��4	��\����d��DH�c��=�d���I�5�zuO̝ٗ|�%��Mg���G�#G������;	`g��t,K���DV��[e�hmkoU��g|P�R��g���I4�B�h(�6��u��-���2ڇ�p:!��+k�r<�Phh�.�׼,q�r��Lt���]4�	:Y�c�n�͒9��(o���@�A��)�����#t%��,�?��k=`�)�J�S^̀���g/T
~(�ӻK���Ums�̉׆�l��-]���̴���Jô�*��г�j�{�,!�����+��c����#���Ǿ�t���l���!�\Y[��o�n����U�2����!�f�;/�w|��u�c;���"Vw��=�x�s��B���l�AԨ�����9)S^	OjG�31m/�8B��as�'T�*��ϡ�Z�״��'��H���"a|ӏJ�<^)?�~* �l�N�Fz����[Z)"�%� �q�QCp%��s���lZ�&S��n�z�)�5�Y�t�[M'���\�o"om��`�U��Pw��0y}0��� �]!±ٓ�h"��r��P̬ɀ���y�660J�)%n6f���j�y6u~:�h^DP:�{z��4�7xZ ���dߘ6��	_��l˟!>�)�#vJ��h��26�k�D� ��O1�V*2��FO�Y��7֧�Aк���Kؚ<�T��2kK6��2XRB�r*%�UB�_e��
������Ӧ3���z�a��g�웒BЃ�/�M1��P��58�t�@�,�V=QKn�@[�i�r�vc��ڸ���5�\;�w�_`&;S܎/�x��D �+��4��L�y�1��[~&1��-�e�f�W�Sg����:لd�i��d6��C<D�\{ _�Y(������ҕ�n���L�V����M��8�MQ�wf�VL�dG��ׅ�ƴ�g,�/z�l�Q���פ
қ̀b�):TƩ��*�� ��ի����E��	�y3�sFϤ�H�Q��O�"�h�@.�G�����Y�
1�^�GQ#��s �@7M�wU��l_3�`�p�+���z+C|��N�3�nv ��	_HS;�|}��7�q�+�����I��
2�چ������b`
y�[����B�tpQ/y�_��.qn�n�$u�V��Y�wG�U�9��Sxj�����L� �>�
�/=��r���b/��K��J�>�� �#h�􆈺�)"�R쑨~@�d�ovaX�礵U��������*��tUH0z��!���g
�%���4���/0�&K}�d9?�*azfќ��P94�V��A+m��O�e�i���g����>�s�A/p��K��YK tgj��!�T�2M2�vω��WB�_���ν�
�F���mgZ��!,%Wn�yD��e�;����@ԩ����߻�4_
,���JN9������֧�a�`KbR/V��.6��-@ڊI�'ߓ���~@���}�5���R�	F#wN>p����
G[4tk�m�q|��e0����l�ثy�1D���/�R�נ�a�Ӣ����!�*�����K��2�����5�c�GP����h#0����<��!�ŔV���lV��0�3��@a�����))�v�j~}<S\јn�;�����R ������bN�77<�6I��=�dF�KU�7���Ŀζ�8z�sV ���Ջ�Ր1�[s�s�^�F� $)�'����~@

g��뇝x\���-��b1���P-r��N�R�G]�Si0�zx!�\62FZ��#0�Vk���q�=܀�Q_���f������3n���r�ߺ	D�* ��ݙ��aˀ�1��ʭ��@N��] ū����7��sh�ղ�"n��|g�'���f3��U����/y��*�0;=m�0�|s}.'t���e1o�E�灤g{24��{��w�Oomb��6�؄o��Њr@/ȗ��u7EMO���^	���/P��x]8%��N�
`'�Vp"xꩶ�@_5D�����Կ᧯d0���0�\��_��2��,~���V(�))>N�7�Dl��#�g�:�;�xQ�4�S��L��
m�և����aU�l�#Jv�'��>9U ����������ܯ��� ��wW-����q�� ��ל~�)��
�WxT�״�O5ؐ��Ry�e�B����]8�E8Bp����Ϥ:!*��AuB��vk�4��%��U0%�3�F�y���*�S"�n�Q^: %XZ����l�˪��jm�y2�NLH�>����ږXga��L���
��~.��X��u��k�"j:r��ƨ|a���x��:��E쒝� 9�}~3΂���;Dc�%��z,���!�ni���0<��{�?�4+��.�I幬�-�@>7�����|x�,��s�`�Y���̌�h�r���O7��)����=j�����P�]l���߫򜳕�p6N�q"hyJ��ȸ0}u��}>Xf3��t]��\ah�9���	ht!`
g��IL��%�Wy9�8��/��<�䄅~f��i�'�8+�Nʷ���Sh�3��,S�S#�L5f�@�d�9T�� ^%z�N��O(g�L��4�Q�ل�t_����"�ڗ7����.:"���S�����+�zV��������%��
��Ȼ[QA>�i�1I�M\��ut[!N�m��^�`/�Y�TUR��f���2D��_*�o�l�1�h;��_?���J����[���+�]�`!k��vv�DZ��J�"sT��M�y4��rOC��h����KF�aP\t�`ҽ�SFr	�!&��Еz��FC�э�.���eÙE�Y���U�"E���r�>��y�bP�c�}�g�T$8�I'�m�q.Y������ݟe��
��/��4����5T��;���Pl�����s�I�qA'?�4p�KN�s��q�Xz[�J�4�K�5X�˷)����Z���p,��Ѥ:<�S�K���Jk��Y�nA\BK�O�@$���Q���2��Zu^��U�Sy[�=�#�&sM��"5ߏĮJ��U��zE��L��r���nb= �J`�Cs��%�d5$/^?���H��X1������co�� (H���9�Ո�gC�b��x��4��{+p���(|�pXd���1W�7N��5s��|j��d��=&�i=X��F/[�r:(�G���u�m����u�ٕ�aǖ	��x��EA1�d���u�:/�\���9��������Xp7P	���	���{�b��q@���&0���a���-�3��N3��O3gG�
?���� vNz�ƫUx$6&]�[�v��\6g��V�]�G�Nl��nl�)V�>V8��}jd�8�޶��l�z��i?If�F0�̈́ǧ�	P������p�62W�Q��K��P=;�(9G7ŷa�f��0e7p��E�K�"�`ػm��<u���Fl�3c��;<o�Ȃ������A+�p\A��1C��(�!d���1�J�BK��:�Q�U���E�0o��H`͢�������x�*l�5ِ�i�N&��I<.��LP�&�ݬN|t�^ λ�o����ы���a*�E���Vnw>Nq�Y�\���<l\&�h�(�'�)$0����^m��>�6�Iԏ+h ��%���H��j�s(`�ʓ�rf��CM��!`23H"�a@+'�0)	�J��58�_��Q�=�/��H�/�^%��W�gtjR��9�Le3�iT��d`�M���$��j}p���Z$�o��U0�KӅ�"-��4%J	_��@�
�9�TO�ĉR�y�f7�Z�f.��h���<���G1�v��S�����V��-��UĬ��n�y�.��^&�.]�߱B�������7p�Pi��>��`��<a+V�Zֿ|�]�K��'���7��Kg���K[��V9A������K�L�SW|�le��Q�*���G��c��NW2��H���H�5_��>�l����H�?4��(lZuN��o��h�F��v"$��o�:��h��5�- ������[��迹��>
�h���Hqw;?8���p߳6����	��#�?Ry������i`�2MWQ$��2��{��H��3�b{���L��Q��_J1����^����c�]��ݨ�y��{��q�O9���sv��Da����b\�A�2���6Bi[FN.��t�&.��%�b�u)g��l:@ݏ��*�3sh�F���yk��w�Aj����#�ba�A+&�oǀ}�ꝲ$�KJ^8εb̅qt�Z�,H ��a�u�Ye������<��o�,ӂ��T�9hL�H�=h�ב�P��!�M��Ʊ�#���⛱ԯ�����ʿ9��sTC�'��
R�|a�r³ϔޒ�Tٿ�9A� �>��/)�^s�h)"�@���q`l$��po챈n�T��7��O���9S�\m��"ZɑÙ��n�S�<Q�W�kH���E��vI) �>��Y��V��&��J���\W`���:b��~]/ߡu����X�M	��h$~�GBhQ8{�j�������(*z�ݜ{��3%R��]7�o��������J̤�蝻22�si��x}��5�8������<j�w�%k��
���As^�qa�QŠ�O�C�J$5wA����<m$��5�X���Z!��E�C����qG��������c^�Ϣ���AMX�� �n������CQu6���	��0)^��,}J	��htW0[]Jlb_ ��t�#��r)�a��p<�����S��@�֌3���k �+$d#|k�f���_t�Ӧ<��*4آ���Y���V����Cܼ^��]�:�Ȕ��;Zg�w���N]�@SP �p��ٲ�FB���n�V;OX�_$�g2H����Q`�6t��B�i�� I���Ak�o h�W6�q�;N	�5E�DV:�pV��e�T��5��Y<�5�F��	׏L{��
������=���"�H��d��G;i��
Ճ�-����5ٓ�亳�[�?f��ϝ &������)n��G:���
�0i���I��X��)�I\�����:S�?���s�~��a�%�\�%Yv�q�� ��Ir;W�V��������SNC�w
k�R�F�
����D�
s��.�������5+/l�Z<�2���T�����פL�k�d,(4������`C1��m��3��8ӣ��'�j��}9)����2倴Gq�����ed�⒉� ��4�r���솴���WMD���J����^��ņ�B�+j�b��j��ǬX#�݈̹�Jʛ��1�o����x��Pn�Bm���cBmY�� s�AВ���z��t��mN��%��&�g�W�B�#���?y
!�*�!�ۤN��C<�p�@v"�ÿ�X~*`�X����L�O`8��W�<���MA6�� n,%GK�K�>��BM����I�A���-c>�_ޛ6`�(����e��^���8o��ܗ�Q�j$~�ݛ����ع�O���ER`ԩ����q��dv'I�D�\������qW��=��(�+<��S�	j��o�X�>�,b�	��l�"�9Z��WH���������X�j��c��YT��A�DbCjh�&pɧo	�hw���Gf��U
9A��'�	A��F�J�����\��3�!�z�B�,*���J��g#D/t�1gS��G#��Y�B����0=�6O�����k��ϸF�Lz�^.q��u���s�����6�@#�r�+���7+ZP�G��GDX�S��g
����� ��t<QU	��	�x���2n���Mr�ϩu�$60��oR�g����������Q@8״�Ʊ8�iLZ�%T��L����b�P���C~/�¯iԠj*��6zĸ�\ay�	�U����wK/�0���f�.�2qL�V|�g9�����	"e���$�+��h"�p��0t�g�ډ/�y���SU�o���$J��kj�Y�K7�c�jͧ��̥�����m�x�W��D<�--L~���a���6]�%�g����g!ِs�X~T�����pQ��Ϧ�=X�NU���੮Dw�[�.0�k�T�LA������sOå<:�Y����߁��<��iL^֟�U��Y��q�j������Z���%u9�p����_$]On@�i;�lF��NۼT3j�*!�Q���]������VhA ?�oY"�n��m������8�bpVY[��t����p��9�=�S�ԧ�w���%ܒ��_��	���'�6h�^���t�6�%<WZ`~��d�I��h`��*�ne#�_6Н�b6�p���N�1�T�H4^v�y9�?h��	u{L�Zo�9z��̎�%���cD�����X�����R3��g�M*دYs7�8�����y���z�iN%�dr����`����6�E/�1fp��
��C����Av�_�G�T9Q��1�����~�9��ScaO��|?D�ΟN6.L�H:����J�&?}��q6�!r�G��4�G0Պj㸜�W�y�ɌsU�C����g�����^H	�A
s��n�_)ۈp>m0��Aj��F��k�I���I,�f������>,1�c���E�O�\��yփC���-����6���G��"E��;� ���dr9
�W��|swnKs�Lu�=���ӟ#$Ղ�|(�6���=b5�#�)j��;xj9��;)�
��g���ZB����g�Ng!V�ҋ:蛱��B~b:� �$`n�@@��Nw�m�4{��Њ���ر���Z�s3Z�C	�����2J2PK�t��]Ӻl:�e��B��/��6�+a��~�Ma�G_�?��uZ( w=gg������tL幤e�J䟸W�Q&K?�[�_��/� b��V6�'#��:5s�P�ԪP�J�Wt+�	D*����0�g������ƻ��̵���~qL���d-�x7�X�ȏ��N��(�h�P9A"v�d�s�V�dБ��o&��+���G����D8}X�r���oZ3����X��h�g]�bܻ�+(��pћ����F�e�V@5���Ed����ۢA;�	�m~����=�����X�=�����W�/./4Q�t�ZՃ%Xib1�/�!|��S��~�f�@�Cji�GP����ϔ��������{��C�m5�Vc��NE��Iũ,0&���?5��;���"�T�J,5�KENQwަ�mA��g���!'���5��ż��D�ژM��h���Ŀ�(�����\�~��]��~���4e����g�0@��0J.#�v*��j>ݽvh���V��4�<}3E܏�U\�o��p塥jo�%]i���A�&O�$i���m���,���i	�2��g� �_B�a֡oۄѵUѪ��ff	�SH�0i��m����Fdb�:��j�+�ҾA�&A��"��*�.<ݫ��5��,��YϤ���E���Kj��J��܉	�QQ��r3�Fd�^��5�]��}Ȕ�	E��K��s>�]�G���܊Ү����1�����sہ�e�Tl��y�?���g!���T��蛙NE\�2� ��!�!`E�;��2�Zv��+�kO�S��D�6V)\� Y��۬w�m�� �@�|965��m�)�W����@!`����GA�+��W:�$��C-?��@��"e�߽�����*�-�|�Uoz�L���K-.բH`�V%u���bz+Y<��Gz����&j�F���3F7������!0e�'��۽����8���h(@r������%;MKA�Q�'`���'����q<R7J�G%+��/�H��x��Bjt��<bu��!س�{E%T�k�d�xh,��������ǘ Q;�<��J�i�.�#�m��gM���#e"�Hx��i}�1�T��G�?�>�[k��B�}����z'l*�p94�YU'�9e!��fβKT��� ��;�N�?���=DXSDp��­�Ru!?I�<<(<4�i+]��6 �hIGՕ����Z��C�6F�<�b��'r�z�S�ft�0�[���ddC�2�ב����|� 6젂��4
s��YH�m;��~�|KZ��n�՜-���U1����+׎N�'�\�"��#�g{�U�*
�����
��{a�-��x�N�h�u6G�"��YYx��?2��ŵ��gX���pSX�s �O�L&�q��-�e�>'�3�v�
��~���<��ԣm��Mk��+T���a������w�����D3a��%L�;�G´P��0�+$N#���Y�->��_q}LÉ#�1�������������!w�Kո��t�����dD���2�rn�3)��l���t��L�q{�ȣd/t�P?���#�uա!��Rҿ�^��W5�
���]s˵�E�ir��t���� s��"B���&	*L7\<��"�6zU�rg�l��)Rn"޲Q/99�Q�{�f/*a��]������<<mpB�
�XV��@\�-G���;Vd���P0�,A583���h�����Q$�U_�د� �R�d'Y�\ �7}d��V�?d����F���� ���� ���)[ ��T(tX�$��'{�&c$hےC e����YBR�1@���7�ԕ+�{х�����<��#�����/N�{(}��^&H��EP;;W�Vh-�o����tO��m�8u��԰��ny(߬�s��3G��1qP��0���a�|����J����An�vU+r\pxv79C��Sxj��ڻ���#*�&��^]*<l��i>�Ӫ�~Q�fv/�o�/E�jp����0x��O؂_Ʊ)W�)����v�&�d�����<k��L],l����>-�33�a�-�{�v�r>��^]�J���o����*���.�h�jT#���(�9$�r �W]j%XM��pw���o{���u��XD/]��K/)�-�o�����5��x֪�j��X�1��b�]����2��SR�zҦT�[�[g;1�W����͉�eGdH��g�cJN�m�-�1�9Qq�1tS�jWe���@�u/��j^�}	>#�<��a�]_��� _ӜF<|"��"�^�x��ΤM��%��̩:@$��}�� ���v&^��pYQ��� Z���I��}j�r_Z�=�mk�mV���|F�s��{<�c��n���h�X�'0�$V��S3���_���wS��̅�	ĪØJ��,Q?j��?�����ֽ�ዹ�W}hVSQFc������l`�b�h��A:����I�h\���1գ��ns�;���C��b1e׭��%Li���ڽn��- ub[k� ���{���d�T�X�$)G������69��]��4�e��N��$��Q�R+%�{G���:�M�v���� �o��E�_��(� t�9Ś�Z�P��!�T����D�J��5�Ć�R�7��+wt�p�^��{14Gf�N�ETl��s�F��( ��b�f�_^y�9H����ɭG��s��ق,�]��7��Og���,#���Iv^�h�O�t�̔t�	L�[�B�|�
A��!s��]i�e���E����yh�9�I�+ ��}���&9[vk��c}��j�K�,}�����	�7�[��1Sl�����d�����6'��L��}I{�eM��a��V��T{X}7S4R���'��Z�l�1��v��?e�jy{C�%�#oٺj�9R)c���Z�T�~�l;�0Re����ro�k6Ofgq�&���yS���"r��] -����aE	��̫h=��x����8�8��㵙��/�λ1�ڝy����[K�Ϩ��cxj�+��܉UC��ybz������H.���tyʉ��+/O.F�f�۬����믭�'ׅe��"�nQ\f�u��+(���n���	㹗�F���N0gg��L���V��d{�j��r��}�¦K ����K	�/�`���'�>L���sYd}��fƘ��3�k8��p;5�o�$	�k_:+T�\b����%>���ˎ�9ð��.Y�	 3�I�1�%��D�������Iڟ�&So.�3�RiW��ק�e)�xw
-1�"A����S)��������5r&��"l�a�aOk������G��^g���3LH�`�7�Uʂ��ưzݐw�o�H������l�����8�$#n�����ɯ�u��4���s�����Ӊ�A-Ǫ�V,������f�v�Nfg>U�+�'o�z�{�˪(�M0bi�����|�C�d��.( �a .�=f���^�I��T	^��ܭ����y:'�g��Ծ��vX�������/4=�,J&�]>�q���
���n#��z�!$�|^���*��
� ����7�Q�*ur��ALÕ&B�h�&�������7��'!�>_�?����)�=��,� ���bQZ�Hv4N8E��7������W�/���tZ��^�n��j��Rt�Ɣ-�ڪ2pL��y�4�À�?�ȪYl<L�j���]>�����UUx9�x�&�?X���^&�j�_XK�1�, �v�xG3r�%��nhj�"o�WK�5�mD�贩(kX�#/
yQ�7�U#��{�o�P�tA�]��z��K�ZNݣj�Q��M^�l�ʨ�'��P���l���APC�"Ẃ���lw]����ڞ6���a�g+'��1�<y��:1Lg��w����׽�^�V�Ҝ��vhΐ����z �6�L~��Z�E��뇎�m�t_#����ک�c���j,�>@������`��� У;7�2��!a%ô��5�(�y�������/�SNr��Uq@��n�5��	G�?�O���u\z�Ҋ�a�
u<�� ۜp�-{{o��y���r��p��:ao�K_�.	�ԏm�Av&~���l�I�l|�)� ޝf�\�`�����z����p��L%&�a*�������m�����`M��;Ċ�ӣ(\qC���h:��Tn%#-��d��U!=�bаGy�'>��B�Y���4@Y)2ff@^�$�Ti��v��,��}��ң���g�C/��5�:ۡ�׎��N�(8���hO�����j�WzR�q�3٭N6�j�:ٺ�����K ���
�z�f�.vr*�W�Odp�q�x�p(��{/P�T�I���_��������g��jJF�D��ݼ��(��փ7?���䏲i,���:4R�>���������}(�(8F�9�o���]�P�ꂳ݌���ujL������U�B�E@1�9����!��G~�� /��3d잖˷�\{�@��p#8��&e�� �� �^���3[��=ˠF��üm�;�n��c�/�$�Z����y�&��D��C����R�-Ja�F�ތ��84��Y�[�������[��7�F]�2�rM�`_�b��!u)�q�]�����ݾp�<:�<�)=��F���O��j���s`W#�}�o���u}'{ej�ɰQ!���
V�@E��l�D+���x��v �&ӇetjR��<3YI�'33�F[�9P�V�{��b�b� \ 6�m��M�$�FsEh�]4
�kJ�*��iD�-r�j�`�K����(典�=� CK�sJ)(7�c��T�p_���v����rе]����+d����rU�݁f���Ň���H���v�O"p��3.Dz�_�?�LM�z�8v���Y:�$5���C�7Fg��9���Ŭ'��v��2��F��8|���ni�ͫb8&�2
$���n��V��
����`ۃɐ���k�]T;�^Ew�D�)l�B�Μe}Ő�ʕچŔr���n�4Ԕ����(&lv\ξ!�<\�8�D�Bb���&�������!4{t�\�4o���r��J�:��i44أl���L�mj���*�vɜ�C��E{�) &sg"{ۯ��+32�y(���~r�hnf�d'˽�/��P��},��y)�s�\dR�$퀾D��W���MM��� �k芪��0b�H*�4Xr��A�$���HK�?C��M�e$�S�B�d�z~���K2m{􉜪YՍ��6�	\I�����A��tsw'b� ��#��������Ir��X(�uQL'.Ŧ�R�NQ2P�"0�	�b�>u���\3�b:#I2ad���&�pj�i0~)�85��)lT��XG�.4��)b�l�ޢ��d�MV�4�$�(R����݁tԔR��<� �`���Y���U�L�%�1R|R�?��]7Χ(Ʊ4�r������r�aC���Y��-�Ǥ�t����lv����|ۀ"T��7@/H�'����[N�o��j Pu>E��V��dǉlh3��`,�Rޟ�G�K�q�<�<e^E�2�bLfDY��p%��`#:�7�5iZ�j+#C:��7�\����¢���R�g��3�����T���Aj��><�锓�/�Ҡ����n��K5]iY1�W�$���˖8�EiS#͵�{��is� ��	�,fLZ-rvO!Y�W�����9jk2(�Ӯ��K�h7T��.��RgI%xj�E�!� ~^�@�S���Wr�����?����^�j��&�{A�2�&�[t#IX3��?����l|�؜:�I.�;l���K �q<�poB�� ����t�����q�A��pq�r��jt�&�U��+$A���6�/�V�`�د8d���q�Ċ�r�;�Z�%Ǯ�#��/�=���4Y�]V�>J�儴�9��^���,(��u��0��UZ�b�|��!P=yF��~�-1�ga�͚c��O���^��aȥ�ބĺh�PE3�=C��K �r����[��ߣ�y��¢�ޓ3?�W��u�x�U�ȏtu#�������K?DƼq���� �e���:e2�t=� w�n^˱����F�dp�O��ڭU>�<�~�&�P�����E_�8q.�C~��n��w̖y>r'�O�<���y�X��pl��+S*��0��[>w&`7�y���-|U_� z��xT&C��I����g���� �AsI\V/.|@E^��\��6�q�-[C�dGEEe�	]i%�`�-��.�>m]�0�O�Q�l���ʄ�*�� �z��?l�v��N\5�!F�rB�(x������Sg%oq=^���g���˫��6;`�i�=	p7c[�:��9� .��O)̂+`D��Hb��]��b'6�)`�2�f���p���)���_+2��#��a���4��]f��l�{-��M�u��ݕ7��"�>��+N�	��b�>�*%�P��Hk�_m�Ϟ6k�>���t��@��>���!��k��x�Z�粗U:�����l�%����w2�� �����~�f/��MH;s�����~��f�۱JUOĐ0���iUT|v��i�ά���,�OGw-jn�t`������@��H��� $^�_H��� �����1�|9���w0�6��{,'8�d��dP��db�RY5�zf�W�����n}�3��g��+�_�Tn\j٣�QZ�^���Z�1�0z׬�[�VYT�pG�o�)���Hك�܆�VH�PǍ��58��Q�iz�	,e��p��H�6���( �x��1;�7 )��d��Q��7��8�$�-u�6q�r6R�l�D�.\�T�����B���ە�-?��D��6�f�=�0R (9$�K�wK�!|K��~�8��«Q3T��=ܓ��&�ui���ϵ��`����Ti��ge��ܾܣ��.��o:N��ۯ@I�1�rUk#���wS��t��7vn�́�˺�h���g���7���}Ic�7g���1���P3u}4��nQ�ߊ��!ۂ�G�Y�!FJ%�.�xr!���(ݽH�eo?q~�~/���_�!��ҫ��H��9FwL*S�J5�K���I,g��`�bf͋K�$>��3o����L�f9�5�(! j#R�{�����L���Rk�:%�\^%XN�g�A�<��'�A�n:��\��a|� �c��7l�<
Zm.pBi���e�2<&:7���ċ4���ڦ�:&iW�[����&�+����{�-�?�
�WO��"r�'�F�K>P�$H�p�w ���:�a�Ά�G]�G�:���,�*�� ��L����/.�;ҝ������(�~��ٓ����Dwl���{�Bc������
�%��������N�v�ݡiخ��|�R���&�p�:�m���~��t�؞�炵�[b�E���\��b�}M���,�[NS�[mӪ(��i���	�>�A ߮��[]յ��:2\\��cy�G���f)!L�Ӽ�B�>U[P
�B�نh�����ޯ���Pn~�2'�q�t0�(���iW���	�!ˍz��J���d���F�d�ԮF�=v**ꎭ2�]0��*�;l�l�  kn9�Z�I��~�;��"���6.뾃f�9k��U����f�&"er���ٸ^JhP���R�͂�M 1[k���w�oz+b�2e�ܝ��bA��%�����b��/&v��;+Tuū�э�-���o��ZJ-�_)Ŭ��
�z�@7D�>i[�����ș-�����r���T��}wV��Ĳ�9�J���e�ٕ�x]�mH�JўO^�kF��1��A��L�i8���"R���\�;eq��fJ \�������Bg��q�Sy�s�ԙDN%��	���b�*�c��{i�oȤ��1���[鞻+�8A�th���{f6ߠ�A�F��2�;b��W�Ԛ��Y��!*Z�[0F��`!wѹ�����n�\^ӝZ�q�%�����J���^z57� �t`��f�c9(�x�a���^����m�3ə !] 8�]{��kBb7�S����X�4~y�5y6	 (�q�w�E��1�E��|Fk�6�	�vÑ�+N,���G
a1�K���V��j��3�?aC�Loz��)umH;�Ub����!<�pJ����{ڧۻ�@C���fMK�;OsQ�=V� y��6�|�%o��zy���;41OL�O^E��p��`�n'�-���|os?��� ,
�[V�i�p��u�&/�����$g%8�1V��:�da$vRY/�-��7��%6�4����֡�>{�PEǫ�#�ߟ� �t�E�$�	��1_�v-�A�lv��Wx�,z��<d���P팲�"�)�=v��ɟ���i�]���������C$���/���#)<�?�1���J�4��q��!(`$��F9����Ds����%�1W_���G�o��?�� ��pA�n������c~��6#�'U�R��� -)�a�k:+�G�w�i5R.+;�f���JI!*�ik������o��AKl[��AHЀ��Q9��8�B=�����#
x$��E+�9�]�����>���օK���*iɻ�w�p��vHLx� ث������Ѐpf�akn��*�\�D�!ѶMI3��i�v������T�V�S�G�2#2��3A�<r�����nB�x�P�$�O�.$��ܖusf3�ΐT%> ��2��lR�)�>���ںcͣi*E�����9YƓH] x�����T"�xYcaØ�>n2�IC�O�L9��Lj;T�el����u*x����8�Kr�ˣ��#��c|,s���	
��w�PK���=}�zN:Vrr�� �ړ/Ɂ&�G�jܑ�b1*K
����C�ϣ��$��z*r����:��yɳ����MC�����#��i3�{4���gK�W4�O�޻|�S��%`"�QsEs}��A�(1�NÔ4S���:r�Y(;��F�*�����S&Љ��W��"����:�/󪹫S��E����#�����M��P�1���N}�/6s��8�T��ѵ��\ ��o4-x0n�"� W���2�Cx�]b���xփV4�
^JP -���ڡ\�h���Np�:����(S��`y<�Sϖ�$0�J�ӥwF�b���4����� �/5�d�"� W���HvW�fU�������4dV�c��-X�غq�@�C;d�=��>3��?��4�i�i#�+�hoq��X_9<����ajv��D֠-��G+x�6	���=�WN�;��
+˞kD�N����s���`Ĕ�¯=8��Ȫ`�p!�$?�[S��-��"�;��$�eȍg��_Íǔ��u/JP�����:nGg�aҝ�z�|�l���c�U�1�7���KY�Q��IgC�=ף�`�Ƹը�b`'t�-��!����Ͷݭ��Վ�!��93Dl�K����Ɖ7�?�q�1��`E�����a����>�2����\;I�� �%Tn`_��4ba!535*$���	��%�7dqX,i�������l�n �T�曠�V�����[��S_����'�D�0�����*yd�B���Ǟ�l�۪�-:����;�O�]�?�UO�Ѧ�f~�=�k*��R�0&{-	�� �_�,>�|���e�$0�ۼ�6s�I���a-��mp��s&0���P��`�G������I����f󊼫��m��u��I����;�sF�Þvk������̀>�BPۥ�mA���nd)3I��2�ܔ�Fk
z~�Y��v�hX�%r��yw��R���~��&�
ɛo�\@�C�z�)�������ٶ�N���Jo�`�����+T^�=��g]�spݴȨ0�ڍ�=����t�!�Lø�d��8��R�oU!��#͘��hg-��/�����_����y$>�-j��+Z�+���Y:Q���q�ౣ�Z��r�q�zY��g-?�,�;>U#�"+�7y	&�+�x�����M�_C#���"Pz,���cZw��&a�j���><�����mZb~nq�O���<�]
/吹��g��A���P���)/���Ep�����Jꘫ)(����SN�P�j�>�X��fk���L���gYm�z�y{�6���cM�۳�1t���Ҵ��l�`o������{��"��b��U^�EA�}�e[�D��M�X��O�c�(��P���2\�3& �8H3r�c]����q�XxH�)/SJ�Bv�u;7�=-�3?\����@�\C�"�AH�:H֠��*}����E���)1a�o�r}(j�f�sfy�p��%R7��q�seb�#M�}��"�M뛴��c(������9"�|��/�����\�7P<�".�Q��Z/"� ,5��k7��f�����c��UB��J�k߈H;�y��]���Oqc�R�y�Mv]m��T������$��d�T���Y9r�SVZxԈ�r�6zu�^l7�M��3�|#�{+A֦�4C����UB�c� m0~3��j7N���=�NS�!�!{�b}y95�a<[�n�/�9A��x�|���̎�R������x>�'��Oh'�w,!j���B�ULd}�O�s�ͩ�����1l��z��n����/��4�x��d�'��1���a��Db�r��3]'��V6�)e�&T3��F��+�"D\�3�8c�cO������m-'���؀�$�n<Kt���#Tc��;p4����yo�&ܛ�"�z]�yy��f_���F*�4d��~�f-�V�p �{^�"w��2�o6�p�R!ci���;K�s(`� C MO�l�Z�#h���!N$�xk��` ����_I�<qS���KWX���[�/W��$�QI�e�b�r.� �,���D�Mv�Rq��{�L�����\������+����Z�Ϲ���	n�W PAe�}]S7N�����D���0�	I�����Q��b��벝r����T��ô7A]�8=)�w�՛�ne
Ԩ0?Z^�����Z�N�V�U���'�N�_�.ԕ;�Pr=����H�C����wc��Qu�a=�$'B��+Ö���Vļ�ȶ��b-�K��
�ap�RSE O��x��0��y#����wp�cn�a���VE��Hm��D8A��%4Jџ�)d�C������;(ր���8�3�]�+Q�;��i�ʹM��<1�U1�e��d�ɝ�)E�U?�]8$���
��P��4l0j�	~S%�����h����4����Cӗ/9���tg�v�u9�t��	lQ�/��<N���0�A�F��/��/g�ܺ�<%�f���	�_�"N�]�R߄T��-�>�&��{�zB�E�������=��?��_d'#d1h׌z%�D
b�xk�%qF<�����,Mo��\��g�B�ta�kҒ����
eD�0+?;���4ꝲ��y���Ejo�lCX婉�O���Rna�=�Y2�XR��.h [U_�K�����z��E[�t�#<�2�ϣ���2�aB� �>��:gW�`1�!:A��8d�@���2�!�ѱ����$�`��m_�M���1��ZL�w�]h�8�;��߅����o�G㎜a+�д+2��KJ	�2�t���)��\r�nh���]v���g�|�U�T9�>�>0�BqZ��%��tx;�#���Y�s�+m�ֺ��94���D�&�\(#�N��V���M���xh��z
|�$EUE�1Vw(��?�YȮ��J�s�Isdٓ����e���Yຽ�zL;�;)H/&'c~I� �h��rŞ|����iF�٘2����WLL�Z��xU!�A,����ȒOFA�y�MB`u�����GKQ��׵o�#�sC��@�	�J��u{�L��$1�*���|����#a�r������ �7fW��$����n���[�:���`�c��u��$��}��\�JD�>�G�
eb.	R����vo�4�r��n��	tL
K�����!���vu�c���M-�>:�i��h�K���B:��3��,��@���#�XFOl��u����2��*�DGLplSz���V>*�*~�������ʯΙ�`L��p�z
��D�Vےr)!j�~vi�+���C�/S��}���p�ޗkH�A�*2:�m�S��{g�ݼ�A�]��ʇ{��@��,X�So%j � �������}�w9��'d򜳂"�ERޏw*�=�k�%�D@�-�G_�cÉ#�j'�~H^����D(�'j{����+�p�H��S�%�}�<�c�lL�\��x��ޖ�߁֨MKnGvG�q&�:jo�7�a��L���c?��>ا���f1e�>��ct����lHyJ�EM�] ��p��:����(��!V�3����t���aғ�/��k��0���&�~��A> �Bw�LN&d�;c�x�������Ѥ���2g�˪�%�~�A)_}�3(��pz��"�}��$B��n]�ਚ����}��{�b��%P�2 �o��VN�������aYG�0�%.g?���<��� �O���w�:�HI5 C	,`GL�L=ZY�C!��0xn ���U�|;/�K���,Vp�O���}䆭K1_�
�rL]Q��v��F��\����lRR����[�D�1|�_0��BOV���$�p��T����n,�5`7h�Yx�-�' ���	�|�M���݇=�.D:�j��>o.8��ϴg�:�!E< ��>�Y���NM�"NqV)[\X�*0F�&*�*���w#�!�$�T�H\D+�d�2>O�P�U/�c�K�?��[+��W�:���'��s��E�\��� �iR�lH��]�=����5dnB�{�P�O��_���UE��0*���q�:I�m�T+�\�@�J�6@�#�f�,h�ᖭV�1���0��_��N3����kѯ� ��y�pk��ϕ Qx�r�;&��)��K�ic�>�/���a쳓b@W6f����g?�!1]�$9Ԇ=���13��9#f��D��x�8�����B5�Pd�R���h��ޫJ�uq��6��4!;W/k*���E2i�anrM���wإ���\�鳤�����Я-����#�Q&�;��y;e������pu����ض��}�<��T����klHP�;�O�YdMhΈUFJ�U2�tD��K�Q�7jA��Zl�Ư�'(�� �9��u�(Tص9�D0²�~��w�$2"�˂�W�C�(L�,w@j)����}FԜ?+���`�%޿��Cp�`���E�tD�@��~���x�m���:�'=�`Lc���;�[��$�	�7�;�\��϶��RP����鎴�a���gglv��@���-!���.�ٮ���5���#�ߛI�h�4_|���Uv�<N7�P�+V�P	�8hϾp������ \Rs?[��ܝ�����é�����嶗k��k�c�hr�X���x"@�t&kʅ�t�|�-�r�u�6N�-ɇ¥��ǝ��X��R�/�]z#9A���1������i���{�
J(OYY0���>�<���:^���AO� ~����ߜp\���zv<��f�5Q@� j�����z��9	�`��3�bb���>����T2�^6����0��Pר������R������,ٶ�w�s��)ӄa>�1sh�d�į��Y��VV1� L��qj� �K	3�ޮ�.�B��rX�wE�5ҫ��*���p������.�P����K�&���m�:�:����Z�7���]m�_�/����/$���q�5+���(�k<�$��ý^<%�ӆ����}��wmPcTfD�B-u����tہ�ܹv� ���]�R��jKvV^���
��v������������r���`�3�����Q����ʟ�3.}c4�)�˵��nz\�`���2�u�'#�S%�c�ۥVh"a�J��ڷq������Z��/[�A����K���f�F�,��=�������Д��D�'�P���⢓���T��"W,u+8&-��H��ɥ� V��D)H�i��͎{��id�� w��թr}
�y�~ԹT��%��@Z��(����{x��\��|����b-������H�b�H���И� '�@� 4�d�l�i�����T�ι�I�Nך��U��&��Uи��J��vt�!/U�-��r ��~N�W,L��4��Z`a  ��t���v5ϕ�G�F0N��e��ur�&A��Ϯ�����,�
.T����
���8G����ʤI�Zz�s�%�_�~?�qb���Z��*GT.(��*����AX *�t9g�����l�ĵ��T����,<�u��˄�����q�;���Eʦ�f�6�<��;�`߭@�n��E��<{�2bTԽ��CNJ`7\�Ժ�>�D�[w�	.&vzД1�")�ŏ�SXb����8��upOd�`)�����.��/�G�����}������Hl c�;
?[��T�p�ؿ�g��F�-���q�Qv
�J�ˬ䛖�Ծ�,�w:�JYh�(�U�ga�R��z�~K@e�a���-�Ƒ�0�k�2]j��Apv;,��̴�|}�3C`S�����t=��b!���~iZ����b�d���O��8vU>�+��o.Z�T�ܣ��W�-�nj��=����߈i�<P�c)~��i��rz���j��{��bAb0����cE��2��m�tP��0 >7�����$���<#��8� q�w�{�<sklO�{5C�AL��������K?���=[g������F8BvԐ����{2�e
��	ow$�ڋg���v�#�W3�v/�*�xWFOY݊��t�^����=�&���ӗ[H�dT��7��K�9BQd���8@�;��F�PaΝ�.��9E�w�JIcCt�k1- j �/�<P�h�V ��" T~�'O�A���[��%J�C����7�7��j�ܩ,ę6�3�|a6 �/��J��+v��0�җ�i=�ۆ`��P�뱵L�0hՀ{�F,˼>!�9�.,�ޗ�`�|(���c�N?�2�/t)մL���2MG�4Y��K�Q�}���t��q�y:���B}U`"�y�˨��N�H��lY�*\g���m�I���e~�����_>U����Z،U�:( 09�i�ҥ˖I�o$7�+^փ?�1�[6[�y,���%�����7@�
��pq�qj/E`��Z�cY,�nU�����|"l���j�q9�q��bK�V�k�V�����w��&�b���Z���ne�Ȍ>Ϙ�b�e����Fg��|����k�v�{�|�g��]^#u�w�=�Q��䠇$|�8�D�7�K����,l� �k�E�kT���KB0��*Fi�z�-+cΓ`G��S�(�G�}�y��'ڮ)K�c,��6��[D�/�g��:��i��0�ɧ�����x!�4d��)����l���d�ǠS��,�jtD��
+��
��0#wx3�J�z�wgY#V�����Ks1/�M���=�Z��)0�fI'�5��5����D�
����'�< �UN*7��u�o������3x����}�pB���� Z�0W/:5�d2`Ê�J1�)��o�4��
��
,0yږ:�0�lmށ�i-�����M��lڛ9�pl[()ɐ��ܚ4|�"m�^C�\3�^�dr�?>;�Y��]�`c��������(Ю�	���|�k@�Bs�ic F��Q���U�\"���f���5,A';�;u�`\j���]����h>��8���?<;|np����u S��c\29��~ �E��0[F����Ժ%+0�{3)��7�P��7����ک?r�|�����\���1��l���¿dTҮ�d������.��Q��ބ���{Za�7�2gB��S�4�����Rm��h��X��i���,X	-Io��=(� '�� }�PuN�#@EL��-uچ�2�VM$��bOv_ ��9��f�y�oY��q�/��k��v�hdțU�~R)��B�pg��iż1�^ׂQԼ��YvkI�����ng\:��,b���zΒ�����ҥ�7�Y��H�H6[�)�LT�Q�td��W3�.��FJ�o�qR�O���5kM��}k�a����K�CQ�
������≖��fo)�g�'�����y{�V�4Í+����V8g�]Y��]�*����?��*���:_1DdO��	�k�жhh�.Q3���sx�D7z��'sRY��BD� 8�(5.�Y�3W���6�_ue��_�-�i+���vw(i�`�ʵ��C(◭�g��ZdKUJTpp�|�6d�� �
�f3���=;�;j�XX6؞h���x�qz�����j�y}��g�����pz�F��Z�!g-pO#Ӫ�2rmO ��4��2����*K�B���nc?�~!�ϒG��р�DP��Ɋ��̤34Sh_x��\a�h!X>$����$�[�[GilE���WUU�k�$�����'D��7��d���y]
ٯ�u�Bރ_]���im�r�-#��tN^�$� ��v��ϼ��n$�;UO�W�5$蘓�LX��Z�INNn�3k�K���+�'���fa(zL?��k�Z<�$=�턃��)��ُi���T��K��T#�)D`�3��i�5^?Y�b�i\���@b:���2@�9}:q�����h)������i-�+�d�j�,� �YQ����F��Z��,��#����wkǯ� V;�w-�T#Ֆ RZ\��`��^�+"��k��
�R`~���Ⴡ�a�����w��<��i'�b��8!��mc<��-c{r�� ]j>]6L+ ���6��,d��y���l��@n�Kr���#V�{@1C'�*���* (��Y��Z����<�"�E�����+U�t��V�6���5���Ǟ"��CG�c��LF�G{%C�Ő
#��y�J�TK2H���LB7��N.�;Q���>7�ZK�1��({e�Mހ
e~o&�Ѱ��3&c+�D�M� a7#���Bep�*�C�w�Df���tp:T��Űj$�.���+��[�n���9dh�E{�}�`k1bTdy�6�e��O��e��G�Fl(+�L�n8��/n�:�Av��ۚ�Cˊ��{�q#Gʣ����p�26��C���}/��r%�A?L�r�ud�`����j�-�.��'���36�ic�����{�|,_�5P-NNf�hߔJՌ�M9D�m���%��>_�#�hf.�Z������mn� �4��E��Y��y��cy�d�8IE��Ou�DN�F�����mp?N�������x���-spF'&_����Y5ӂ�p'lG�V7��u`��2�@���u�ۍ��dړv�n˘g�:v.��Ex�,Pݵ�n��U�-��o@1�jy�7��>�����D%|}�:
�fX0^q���(W�_��� �_�����K��	��t��C3fc5n���2{�ߑ���eAw����({��<Zm4�U&�
͜/��C*|��!���-G����ʸa,i(rT��vf����㢜53)ہ��<�Y��N��*��{k�	�~�Ԛ��C�$o'Y�;S�ڮ!�2}�[�a��z���Co�N>^޹z�F���?i)�F�=tV(�}M*������Y2�'|��H��t
�ԍo{����/��N���)]����&���: (���E�b�b��v�O��Va( �#:t^��;�ch1,�w��M���g�ƶ����s3�k��S���e����шP۸4=z���P��ʭ6}I�Z:��h�
�3�<?NQ�2xx�)�'m�5fm�?ƪ��q9�%�2M���`���*
�����8s��m�#�&�0ց��Mٔ�"';|�|b���v�UEX���2���Bd�v�`:�f6a��'��M �ڭ�+����r��F�o�q��B\_5���T�bg�.r���s��[��Q�[j�sU��$�j��A,8�'b�ֶ�(������*���	��`x���,�jM�˼�Y=�P�m!�Xˌ��Bޜl��ŝ�èwĽ�^�G� ���E��O̺u�:�-pk�v�2½��ne6�90��)�_w���X��Ad Ac�Ks��j�7�#�tr����\�O�xξW���#Կ�!Ϳ�J��隨awȂLS]�W"�["�a��K����鲇t�+�#�=& eR����
�5w'Ju��]��I�O�s��Q�ŉ��5p�]w�D�(�kL�@Pf�`�'Ȼ���t5��Ƌ{�\h#=�!�
�kuh�!xzǺOػ�E�M[1�K��?�O�Ï��oG�J �� ��up0E���b���-�w-�������ۖ&3C�*��2��ld�Q����Z�ԩ�ɧܨT 28�y�&(�A|ȣ�W3)@��O2���پ�*���2j��m���Yi�3��!ƞ�q"H���.�6�>�J�~\��Q���q�B!'l��kR�2<7���,�=�/-�������&���2�R���ր�_�+�b&�7P����`,|���^����2@=V�������I_GN��y ⫤/�ȀȤ����e}�>��;:hʤ�Bp~�0�]�M7Y<�M��9�	E�����
�� f*�(����<
2Y)<��@��[d��&�MZ�Sn��eGdQ�V��|�.\�C
+I����s�pn�����V@�.a���_O��ߘ���|�Bwmï�딫h��^*���5J`
�jy_�e&S1$���\S�I��kv3fl�Ν<�H]j���݉S!��OlT*��y�4������?�?�f�����>���q��xV�/��y�~.���٘'�;3d#ɧcӶ,�Zc�����>�Ssw��hF��@�w[L�z4�2��p��W����R\H��r-P����P���d��
zl�E����{R6���U��m�`d�\�W
К�LS<}�e�3lM��&a��u䍎xY��J�׭{n�8����x:���R���M��ZB�lu�a���~B��̩���r��c)~V5WI�����cضQc��:�����	_f�E�g��s� �JoE�P�ҔiŇA5�W���z���4�x�A�)M9��Xn����������������W��9�	P�M��1������X�Г�1��b��t�q\F�i͑���W�ą�C��ns�>:�VLwN]u��9.�K��j~IxE�&Dq�Al1��!9@�RcjH������~A�CY�D�g]�.-���(�J�SG8�N+�2����I��L�&�R)�lc�׳�볭�{%V,3�Z���<1����]X����X�����e�.��P�+�Ɠґ=Ke�z�Ȕ�&v�TS|�Yry
���h%ڬg@������a�G����p��b��y#����<5��V��O<L����=(��4��]�!�4$�N��y.̈Rqg��"3��*�Ѕi��0���zM�	�.Ps���1[�xNC�k_yJ� ��|3��'@�5����Wr�����9©ok��O��@�����boM	`��KvDӂ\Ϝ6`	�| 7�݄�v�a��>҆����x���>�pQ.�+�[�ZI�3l�T����<r���1Z����9�u�ko.I��J��߽g�4w9RT����A��ؒ��]��I����� �����B���2��%P�����2>�����"}ݙ����G��Ӻ�L��|�2�"K4Β7�zR3S�X8�) �Y�-����*��~CH�e+>f�3�G0���%����B�<���`6"�w��G���������N�5�MG˄[Us\HV�R0ʚ2�v�<�xzW
��|o����	���W���퍡,�p�a1׋������Fڔ��ۉZӘ��Dd��D1��n���6�a`�R�~�!�E�͹pǝIy�0��I����D�M����^[:<��1E8���j�a��.Q�����.N�n�k�3���(,�8W�q2[S����䙸��S�^�]q :��%���62
�Ao���Ѫ�"���2��m�^z��v'��5Ne"X��j�Z?� �����˾�Pn�q~�/�M�|���DZ<&�s�qݠSp6,�"{2=��w�dO P{�����>���ԍԒhK��É��:���߸�^�
r���c"�^dPc�u�-��4_���r_��D�YaC�Ahe��TAȄ&�fp�hi��>�X��'�j k|�ā�6�ྨl����bTLȂ#a	���z�r~D�������%~���A��.�_��k
�B�	���O'�I��h��wr� ���5��ZRX�f�\]�(��DR�y�dg�Q	N�CR�5��l��3��o}�{RWe���>�_�� ۿ`�P*g�W��<����x���$�i�4%��(g����L;�w�t�t(�]�nhܙ�B�1�-z�fQ��6����<:��*3q:�ŞP��T�����s�KL�J߿����r��3[����/�xI�i�l��"�2^_{�\K~�	��e�):���O���R4=۟���u:=A�j���$��ʵa�kJ��qɏ�O��')�oj\ ��@�z��s�Ƀ�fȮj%�v����ϘDD�93̪��nh�ppX�\�2�1��.i�}��8U3��̈́q�o�2���-'���75pλ)�H��`Y]*�x7�׽Ժ���j�RΤ(���!�S9:\��$������@w	#�+������E�H��R���E��s/I�'��#��(��U您1��.V��l��U����������&&��xB2l/��m��͸��@:������r���^.ˀ �^5RH�ݲ��T!=#�e��Z��[��b������rR��m�+i��u��qF�"���	��'�OӪ'��A�C��J@�E�pr��tp�ҪH&f$��G�����<\�* ��"�+k��
6]\3;�[D9�D�?�[U�3��t9=�uG�8�g�(��	���.j����Q@�A�rX#q���E�p#-5r&���R`pOu-49=`�p�<P2N��FA�9�`��s�}�����{�lW�(k���P_��d�ܢ�Q�zQ�w�qy>���6�MT}��u���}b�6��k�/�)�K.��rkmjՊ��+�����9�½��틆�+�0����c����m��z�3f���,���&�o���uZY�O��tu@m^)2��X�+k�e��mi��Ya�	A��	̺�>���k������������V3���S�e�N�A��N 	Df�R`�B��ĳ	7��G��P!?]�nf��>0T�mZ�aj2�<��bv���<nG�2]�t��Io��
�س�F�A��ug}�����y-������`h��i/���}m�t$��<����� N\�����X�y�!�Qw��T�~�c�?��gKr��&���W�]�h��*;_����I�J�UN���մK��)�w!q�"!�����[��t�g��DE���Uq"�}��[����n�{��n\L4����`4��r�Xg��D>hv�C�yɑ,U0����r�j:���$�H�g2m����1���*�]�3�{��7�������"�B��b�����[?���$�-x%*\���~�D�%R�����	�R\���])]�z�.%oUG���mCB��!�	��;�e�p6ӧ�P:��]���?~9ȅ�r�� Y�˙�[E0R�Q�`������۩��o�����ŷC���Od%U����*�V3jgq�^���7${tcH�������Gk]s�-�g��Yս��w���٭��|M*w��j�"2]s��96��F<�� ��̣0�1L'��J���#��qg��zM���j�1�� >c��s�=��`Zm�z����y�4C6v�'\x���f���]=ZuE�͜E�%���].��4����\��<�»"J)+�l�i�W��O�w �ߨ����p�.A��(����|�q�9q�%�u�7�Q���1��� �fU�B�m�m�GȺ��a�R���!QT9t慄�+��쌭)����@7;���34��? �Z?�i8�d�֖��`�N�������	I��%,��mÔ�R��OM3�ື"w�d��DA��/�w�FH:S!��׸L���!u�v	�W�}�d�5�m�ʶ]���]F�Ę?�>�7)�BM�8��՞��N��O���P���-�v+kP���t��Z��A��]�
���חy{C�W��MԐ����>�}G� �0c��C2o����x�B����5ȶ@Sم�J��Msayl{?N���2%F�ĢךC.�Qְd��G�����&��:S�t?�%��� n�����1�a�o�n��.��}��:��`wT�X�
��N~n� J*���M����s�\
���g�xl�HYG�	��p?�VݽO7�ġ6P��
��	�Y-�9�_��Cb;�7��MG���Ԟ�A����ZI�F�"$|�@���#��ir�S���Q���ȵ�w�6ɛ�rx��v�ɾtl�K�E�[���f���x%�$;c%,�{w/�L�\/LT�`���+��9	ELs�:��a�&����V1�^dp��!d�Y6��w}1�,n�0�y6檹�W�U�{�i�=��dI竵!�Ct���jڔ���|g�	����u'���}�WZ��� [,���Y�<��&a��:���'��Ƃ�ѩ/�v���zW���5%�O�Qx�zF���2�N�Q�b�6�8�:E(F�h���\+�. (�G׶
"������_ēM5�Z+I��/7U]�C����c��A�yZ��e)�@��>�Z�a�YS��''
��lt������&����Ș,� ��(�L���к�L�W�#8IxI*����J12�X�T�I��Y��i!�mC��lq^"؎�����T������z�邸��B��%��؀�>(u}1HκBSG[��=��8�}��?K�@��v5��O���31��O����
��V�S��@6ǌ���w���5 +���g�`=麲�ת=KM�M�U�{Lk��ɾpO��ZUl��:.�W�y_;l���`kY�,�b�dCOo��鮿6���󾡚��,�a+0��`��ܧ�nJ�܂�ã&��D�m()�N$~d� k����rk�n���}n��(:�sw�$�}?����)o���1Pт�s�5"H��?������7$�����W�z5�Pf�XU�x�M�'l�����`ٟw���B� Q����A��w �n6��c�ǻ�q�#��mW�SW��)V��+XN+�ek�)�n�޴���ƈ�A$׭l	ѵk��n^����:�Q�QI����8���·��(n������?��^�.�ۧD�TU���D?�޿�L/ M�,B{���}���
����Rf0���D�d��y�4	�\~���2�ɸV��{�$(��	^���9���"Ẑ�^�I�Cs�v{�y����ʡ�K�s��,W+��w[��S�t��K����#�.��
�	��s�����1)`�m������Udi�����=����8,|4I��:vM�ށ��8p��t[mo=�k.
kTա8"0m1�u�溠�I���
���q@
'�t�	k��O�lH�m�ÞPH��V}2D�d��M<�5^躩�	��?;�p��G����ǻ��x�)+z��uu��S�����󳵞x���Tf%�D��N0f���,�j39gA<뛲ˏ8L�O�����-p�Ė�ؔ�r�н����˷hfӁ �I����[��G���%�U-40�	\4�`햱���Jx���=u�+��C��;ؘ;/d��3k���O��W���DG�,�X��J����|�F5�O���<���/f�*���>�7�Lq�1[�	���I2@Kv
ku�LU�=g�β~�B2[��mT�Cx����Y����	l8VtT�+[B^��!�ٯ���Ug�\#	@�hex��oѡ� �AD�fUA>o���#�Hk}�w����+z����H�rZ-�pRu]�k�{,�@�Gu�~���^���W,��j���ߙ�`/q�E�=3��DXyMQ��#{��� �Ъ���Qhb��k�By;��l�u��x�a�����2�]|��ݯ�;��ۿ���F����j�%����:��7u�!�0�wT�Fi]ҀϢ���MU��z��R!�D��ܜ�̚aQ��]�@f��F��5�,�l�A��%<��555s�<����A*{`��`179O<"E\qv	�U�=7a�mm(�'Ef8_xy[�Wr���
��s��ݎ�qG�$ �עv�9���\*,�3�8oEʆ^�Q��B�*" ��Q�جp����ֳS���!um��I�0H!�|�	xN���Ma*)���2�K9�?d���N˷�U�c��������2*I�^��n"V�L���_'���L�A\�=���k_��"����݁'|S��M��Uk�Ej;��͵�h8��E��}L�����D*'��	�b�C�	1�H����񫠛��vܿ�P�Oǳ��'�C��O$�YAgsX2�u<L���>:sy��]TQ�G�U�ϲ��x��I�ٞ��(b`��E��R{Vn��:��m�f��ڂ9�q�b�O������7Q�^(ot"�00Q�d�G?�aC�4����h5��d6on�|�"3^�k�$y �q�L!����Ax�A�|o�͘e���w|�i��C����Iws:��=CHQ:\iV��A(w��-.��VS0��? <�Ֆh�l�;��Fϖ�fy�������(�� ��p�Uh�UVݑ��:[=�h�gϨ�O?�^���/%<&�ꑽrj���N�`Zk��A�K��6�nwJH�8���vlg�Nz?��{~z����bw�Aڷ�<|��NF��xm5���
(��^�DT��dΗ���u������>Cࡰ��a�O��� &n�՞+��w�0���� �V���2EG�t0���|1
J|,�2k<�ﰙ�:�(D�6��.�΂Z�:������5����u�໽ lLw�]ԭ�"�����'R����u��X�6�FGE�A�FL��J<s((����#������?yINY�.�w#!n���/vpJHt���R
l	3UZw�9[W��&	��s*�����Fk �С����+u:� ܐ?���3u�rmn'�r�W�p��(�+�п&�,�y��2��u�@�l��4��@����8��%Z�R��U�Z��'�v���)�m�=� -�'��D+�w�tq4}U��:��>��>��P�����%n���96u�,����f��'��# ���J��D`ᶁ�7ύFsճi��E��5֣p!Ȳm����\�z��+Q<�(9�8l��ւ�.Rq��y�K���I���%�f�I�}���,�7�%�"ZK��1[�_/U폽���z��8��	r�P����_�T��t��S� }����e#�����X!f�nd&DR=������A5X��Z]Z�9���l|kp���O�$�^]���B���P�ǧ�%1.���#r�k��u�41q�#��	��ćy(�=\i=��M�í��{]�nq91,��x��+˒��Y�{D��}��8�=V�BׇcBp#���@3Ř�)�6�)dݔ�?�e�<�K��8�rp���'��^��(\]��ǀ���C���$�g�o����*���k�O���y�+)N�\'{�H;H�)4�����YO9C����V	�_:�Q+�\���{(�T�r����5��1hÉmFө�p��_s�֌�2���L�u�3¨�ѓI��Jz�k���[�h	!�ϱKV���m����@^9,�'
�y�sܗ��Aq�
?�H_�o<wE��ز#=-g�?��>�<V����~N�(n'����tP��oy4���p��!���ƀ��t���f�u�*M�џܑ�/��wR�|�u<��Ħ`���b���#پݰ��uT}����|�"�����G�KT������Әm
x^s�K�a�8ـ+#8�Bه?�؜�kL�&�O�"m�Q�u��6���EC�mɖ����V�/� ��Z��;�
C�]u��N�ʖ�N�-����O�9��8g��4���rC ��P��ё�-�����L��e��Ǎvw��#�8����:�q'�Q�ݏ��yԘK�k�~�A�u� P�5����ZZ�K�N铉�P
�M�	*`ͯ�URCJ�Ν�дn�<N�����w�_�jVo��9yr,L�r
稘�#*0?R�
6��Y�5���C
2D��/��d����.ԝXQ��	O�5���L�a�1홶�lnC����~F�~a��2;'g��
�5��SQ6zW ��-�}�kt�F4��񝑿��]�B��i�m[V��#'O�@��j�%8�0@ۈ@��KuX���%<@г�I��rdŰ��D4널�dކ��`�T.,�V0���2� J�(jt`θ�`�]d>���R��EN���O7-�ؙ	�i�u�|�&g �����ׅ�$[�Z6S6���w� �&���%�9��*n}��מ1c�f_u�����J�7�Z������V�%#�LM)R
��S�E/�Nԑ���!�W�O.�W�8�B��V}�U��a9�.Q�\��a2X�1�b������β�l[(ffQ�k���O�J^S�qL�ۨ�c�+}6����?4@*wag�2�����$�}��۩�4�q��!�
�<"�Z8�=bɩ��-ӁE��p���XQ�����A�wwP�KV{�c�c��T��)�$i���@~;D���!��w
�*�2�VY {����I59-�By�������N�ߓ9P�#bu,�:6]�R�W�a_���'2oֻ��u�2�����n��#Z�hC�!�����	�o���SK�g(ß;�iQ�v�Fs_����!�8-\��W���	d�m(���tb�>�I��P�"T���'��S%������z޸<���m���1�a"f*v*h����/]?9�x�8��U�]�īAt4��0�s�ϰ��棋�=|�q��"��ia�y�~����-�0Y�|aw���ߞ��T����u��tk;�j��k�8�֫1��q��ѝ������F2�º���ņ��Ey�v����"F��n�1�$�1�3rN�b��ŜN�6�#Mt;e��QyX�'���T��ۆ�d��m����L�H'F�����bv�C�&�BYKێ�����_�q\�>��G���kPve�ٞ���E��ӥ���Ml��GB�r�����&?'bG���P�Uh|�ް�KI�z"�D��J�S\����TM���B]���Yn��L�f;�~m�����#hl��kj�<f�%��Y߀���T��}��"�{K6�,L�5��,��ũ|Y�b���Q�?���Wǀ�*[˹��ql��x ǁ�����*��u ����R`2"��B�#a�����⑑�*�̒�D00� Kp7B���4jR�H2��Q֓�NXU&ͻO��߅���iB�p(�2�Z��)x��X�5�ݦ��(g�?�P�:�#��r��S�0�����de;����(���0T���H+���m���\C<��.\�U���w8�����$	���I�=�!�Χ��	!�ʺ��5�VU$���=�u8�0�V�%M�..��Q�P��G���m]{+Q\,j����-��E�l���~� �y�]/�9�<�+F��+�)ڒFs��(�	8\ل9�g��`����Ѓϊ�bt�Pd�BN���;9	�':q��@!�c)�;R�`��=��y�,^�b�����T�FxW◍�`*j�YM��n&a �ܞ�t���!�Q�Z��b:������|�e���b׈��=cX��r�������s�F���{�&iqKPt#E�r/gah�^�Pp6L+�@���Y��`�i�'���y��Hi��P��ﴰx�YD�|x7.�;%��5�ϲ�Fγ���|��D�<�#	�Ցx����Ǵ��^n�n4.#���;��t��Fj�F�6箁�i]i籩Bu�U�?����;�@ ��v������#��:#�:Δ>��m��Z0/�.s����U��f�d���^\[{<�B&���L�f��J,\�)�����I��6&0��X�h�7n#0?q=t��f��Ph�Djj�
�}}���Ȏ�SY���.X�@H�&�����9���n�HA�?�\������p��j��I%�.\�^��m����*U�A	�t=��0�}��^T��#���7%�ޖ�>8ֺ)�|�� [���Iv��㟸<N��]"���<s��[	��A�/�%�`��`zT�q�g�]VL\`[��$e#��4�8��'p�N�|r��{K:��k����f	�ғ}��i�Tu�e��f,�"����/�Y ����c\����hވS���,�^�F�w�[���d��M��꽞!eG�rӚF���0���	P�4\]��W���S�6�\N17�O+�1V����E�3����c/�s�%*Ę�3���5��D�;�.�_�p1�5{�p����[|�ŧ��]ѫ3���*��ɓ56�y�/p���ta�����%�͏����"��ӟ�߄%��l��HG��ș�(��v\�1]�W���I��/���J���x0���%Cd�}#�7g�@V��a�@���D��ѪC��@,3�����	�� ����ens�Ф�6�ԋ�X��]�R��n��Yf߷1���p,��Gl�>#����5vVjZ�Z{#)�GÎ�cԀbك��A�
^X��ـD{a�&�xW��F֙�H&������lR���"�B��T���/�J�"��S��2�#@Z���0F�|���f��Fi�-���Ҫ�Ps�ZD�ǐ|���X�����ی�"Jȸ����'��H�Y���1A�p��Eu�I��4��g�n�b�Њ�_wjV>(]7�Q*�I7�����B~��h:+§�F#J��͆�*U� '�`#!m[�	�)�-0	��(�.��Ƽ�ď��w��i�Ove�[��w�B{�d�[l�XR��x�n����|� ���9`ca���k��z��}��6�"�P'�{��(��c�M=�jj���?��4چ�`��z�1�E�~�@�L�g�����@.c�G�yجu�fSj��}ΓC�03aoꥇ�024̷�l��k9��+@�(�m�'5�\p�y�:l�iöi��U2��ˇ���ql�cp�g�Sf�W1Uv����:~62�|wç��^ s�HG&���g��Bo�1N�<,��;<���XŦ��0~7����:wl�F����>�܈�A�|�U�HXC�<qt�a})Yq*Lzzj��uƮ�a�aɎ��ÀUVd"�켷Y�n��n%y������f�]>��;�M���������j~�!��ޙ�w+j�C��B�5��6X��ѥ�c�o�E�t���M2����s_�04;�-rA�"Tr�l~a����o�e��y�hꂶ_�. �9� �ПH�S|��w���e�O'B���!�j��@O"/.���}�}?�V-�j�	 i�����kjWt����\|�$���"�����3�3�U��1ALa��ϖS~�$gе.���98���L;1]��P(B�a,��N��<(@�/q�����"M��#;��r��4���.���U٫���V%$�-���R�F�&nGB������D\x�̐�ĩo�2��|�
Q��+�'�T}��6I�` �����ű�&��,E��"�AQ�"���\����,���((��	�{&�g��|#�~�s��f�KX��oғ�{{��I&ϔ[���`V�<�����Q���Zf8�����>����n,(���&8��g�s� R��22���:\����d����mϮ-ΉF���G� 1����9e}Ob���[�AY�4��hb��lB�dn�v8���3��ozVY�\��iN�2NF_�%b�.��`�F��Ɣ8.� ��ku��듫�c�5�@`��ac��`�Px/3�#���ƨr�O-)gg�u�y�D疏Z��0/͠nhq��c��+Ș~~�e0hLǨ����t��`���?�k� ��6k5�xBYD8I'��O\-��/$��<�c�{�"���e���kLغ,�钦���LI��^]L��
l�����b��6s��r0a��]55��)1�O��0��.,����ܼ�L��T��j�#����Ef �7���J��ДvDA1D�u�q��B�$�X�<����f�烘;��7�?�"q�1�nu�㒡v�u~?4�z'r�+pyy�D����T����muʖD!F�(g��n��r�J;�1I�)47��WDir翓ew�� _�
Bd�v 耽�֜3��,��x�C����dQ�8�5���f}���6� L�A�T}+�V.tѱo�&8qg>�xr�pQ��,c�qt����"�YuW�� sr�k��7�Ww�n����}m�
�a���x�(,���zR�c�L��Ⅹ���d�ߞ��RF��������>vt���K�]<l���s�ά0d{I"z�C�!N�����Jd���T)�u`�)�x��֗e�t�zo�G���1N�V3��!"[���`h�A�p����دD���s��O���ʼG�Y�R&I��%e��(��H|���ZB���%,�:�W��ڥ�9Ƣ}���^Ւ����)�t�W���J,k���>�0[�3xT�߽��,6G�fm�Ԏ����4-A��z����K|�?� �ϷQG�e�
7�JK$R�\ZG��x-}��| ��1�q�dm�S�ew$�T���ep��z}�	� �"�tv"V�f��N7=G��ڋ �e��Љ���޳~Ğm�������j��N�T ;tq�Xp�a�Ν"a�n%��?�lO�Q�T�.ZF�䵕����#�K�\���Y��э�҇;��ě�,Q�2�m�0h��f��{e��0�(��{������p}4�����of&���ω�o�O�Cָ~k-V���>��C!9m-#j�K^"���n!�t�e���NSZ����) i��]��|Ŀ,�<�J9QN�Z�]��\c��ƴ�э�)�$<����?�P��u}=T�|�-Z����^/2�q�F1���H����R�c
`cW�,�d!��!Qݜ����xoUH*�rѻ�GW{"����{q�~.y��=-3l�~|-�ڒ	�[���{�'@/05A� "آ��<A&-��7�/¡jg��hth!����G���\�m�j���56���TG�~{��f�3�����x[��Ɯfh��,�?vB��r��Z�?X�D�X�pz�)����C�;M[�J��ъaf[���ny� ,��M�kAI�`���`WD}|�"����4�n[X|mc��{�D'�.�Pu�ވ����i��޳)�����S�>0��޳I/����Bs�o�nX,9@��>�"��e*~1	��AY�G���o��o�R��2H�,J�!�[�l�H��0����im"^kn��DIg�J����C8{E�g�߶�ӭ.�XH�]eB'I>b�s���fP�h�1���\��hW^��g=���ZDx�x���'`��5�����]  ׍����ѴoOQ}��������ļ\Ί�М���R�my��G*Ƚg�qz�;7}g�f����<�s�{���&��U��,�㵺�!,�a�9#`��CI��AG5���p9n������N���e��.����?	Ȑw/9!�xn� �$�n1Z�M�8�P�s��=��X�\"���	�0�S���{f�G� ����k{֢,�/*%�xS\|���U	@a������lK�m��?F�}$5n�8"�$#����Й�&o(��T����H}�$X�O"���<�~��-����a�~�c������Q`����H�]��&q��(�N�¾�)�<v��;4B�4	��=g��bw�;�ŒB�x<|]�&��aI')1ʻu]u};��p�#�?]�H��W=�C�C:/��xS��&�F�r0UC p�l�~��ˊ������[��4��0{y�ع�`��Ns\ ���c>����	t[X�ۏ�Z�����s�_Oe7l�R2���qO����ݹQ����=�v^�³��ֆ7O��+Ƹ2����M}0���Ӷ*�4��HTT/���h�5Qmd;�����Y;��Wa���b��o�bdD���� �H=Of��r0��g[���ׄ����FZ����*�-77( �*��FSz��/
����J�{~����3��W���\B�N�d�� �mL�YFΒ������*���$鍽=��"�i��b��o��B8d�LT���O�i �����#8Y���,2�ls�~�ܫ/\2�qŧw��}��4@�����UМ@ �.5]&.����{5���~�1�˘H�r��=��tC�+q��BF(;p��ZR�4<�>�T������Y�M��������J�+��� �i@���j��+�b �4�9���H�Cա!�a�sj���]/��P�%2v��W���H�7-�j�Fh��h���%�����슉F���)o��Z�����6�8�p��8��t����1�(eAE�"B�P�q�:Jx���L&z�q4{iř3���m��?v��/�8"�n4�h���L*�䗺���.~�
s�*|:�8��Q���<_L�@n"{���C��P#t�S�xd�2=���q4h��	o�ӑ��L���*.2E�s�B"$ϱBD�-�0�a��A��½�������k�7�Z��{�f>��4��� L������Y���f1��.9{�[�w��w=m�S��ȵ�8 ���0>����GI�*՚qӰ�ӟ�<�!sh�[wv��\�#8�9��O�Bɠ،�	�6;��x������8`�+8�0"2'tK4ZS��֎�J����i�B��|c�f��oU\��
��P��[���=ĭ��~Q2���w1�g1�HL�g�י���i��D��jB�cb�L�*MG�A���@����u���F&���K�<�-Y-`�p��⒓rM?Ċ��/�c"N���8�D�c��j�%�,�7Ae;��a�J�&�I��d�L0�E:�����9A�ҫ�"�a��f`ꜸZ4���'�O(�(TI��7�W�W�Р���ݱ{��<D�$D�u�ɏ`�h��)�YP\M?*��C�Տ���u����N��e�*�9��@��R����uw.��5Q�}^�.����$ ��G�mM?��8h��g�����3qA�n�@И�l������U��2��4`qFϘA��:ig���̫��|���U��i���
�*x�}��~�y£i7� ְQ����4�b~{�CDM)#�]���#N������ �:Y�s��#�ѸKe�Â�6iȩ,	Q2���f�B��	9vqJ�9�8C�D�tK���ln�q!������i���#SNqf��c�b�$�% ��H0#_�n�B�(�D�-Z��y���]tȇ����8��S��Y���3
�7wa�7 喴Fٍ�;�#�]`��jTk�^�[�LcȔ(cj��L��r��_�'X�-@�_��@�#$X�Jz����80Fê�y��1e�-��,X�r�'�4,D�q������-����@}�f�:J�@���:��w�6��w]��Ϩ�s�}�B��R�)S�[N�b�̩�j����~��.VL!.D�N"�@��Y �33��0�	���E���ߵ���1���n@�Ǉ��`C�E�x�����M�p-k�w̩}�����ZO��$�{3�|�l�EDO��I�����X������_#���:H��ɶϬB����g�(+KJ�Y������8������H�R� �08�1�x��߷G�JJ�U$�C[���5?�+H��LO��~Z�#����=�g�LM��Ս;�G?�2�s���v�fL?��q�&*T���lz���qHk����y��e~N��,�t($(���5F�/�����ln�xlw��k�}��n�/�V@��4(�<�&��6^Q!R��3"P�0���8����m��YnQ����,�)�����#�B�)1���;a$�����O���Y��pE|I9+G�g22~=J>-�,�z�=�#�=e#rM>`ͫ�>b��9%sޚ�KEb^�8X��{��=�2p�@ ]�M��#��ؖ����U�vD~vQ4o��O3𵚿ݛ�-�=68��X�&j0��a�Eޜ4��{�-Da��:�5�:��W8nv���f�Z3����7n�����qp�AߵTZ���_��4j�u�z-O�6�*aj�4��&~�|���M�1M�����	�/`��,#%� Y�ܬDtH~���e ��� Hve%s�|Y��N��Kw6�a�i	!Yi��e .��]���	��,��08'������\�D�;M�4���B��t����aVY?9�9Y3�i���@�MD-��\��,�� ���9-��.�;T.uE1��/l����R;�s��:!�}DM���9�?�(��]�6��FbPx�b�v8��6��0�[�R_e��mE"�H�Mv�L��:���:��ɾ���z��;*���F��̝
���� gO��W����|~}��'�$3�	~�~��C��G7�H	c3�������)�-��--։���$��kC,ʴs��q��t�X(��,xS�+�K�����	���j5r�f,^�!�tȊVl1�k�Ҭ�7͖]�����T[g�UN�
TC�u����(N^i�_+��5K��Ь��q�R�*���ӑ]ϱ��� �;��U���5GcG���i!Ilv1BT��
����S2�'W���#�f��L�C�,g}�,��fH������XЎۑ�KD��(s��p�]����>'���Gq\��Tͳ�����#%���9�}���IU�����f(n|n����M'-d�'q.};�ݘHv�k���pf��c��eYr7L�za�:����_~LT�ݽ?9�&dE4�
d?b�gk��ϖ�-=�R��(�������S��:�00v2���!:Ye�J��|�m@��^�s?��eϘl(��:X,_g0��l�j��5��WH{���*	����??W�\��[���i��|���/�nT|GD���m���*�%����2�`4�����+mG[�m1%�j�aw[f;m��2�Ih�&27��O9�[]{*Q83���1�P���%���L��-�T�^v�U��Z���,�����C:��G~F�{z95��R^I�^�⊥����6�"$b�ajR9W�T��
X�l���_�3<��=C'�5s���>L�Q�^YÎ�f����u�	��1ӣ�}o�5KTV�+���'x��z�w��V��o��q-�W��x�s�R�=��\QB  ��z�3)���`��lMWѷ}�8��>�'2�}g�_Ad�i���d����Lٵ�2Bc�n�@�|��bG�7����m�C��E^�����a��C��/_�Y1�8��p�m�h������'˫�ws�8]��,(J�F�{Y�d/Vw9v8�Cg1Z7xk��T�z0>s|5pw`R��E�_��t}�ٿ9����@��jÿq)�������R�nW��K�9�F���04�r��s)>Y�%y�>�W��ҹ'*�2�� PX9|�:�=���m��h��2\ۘ�Z�(D�)��r� 5)r<�׈n� ǭ󾷚��������F�� n9�������g��ya�#w�{^��TjZܛ��q:�ɺo��F��CZ��ؤպ�EP�'hsh��A�f��z��N&�eg�t��`C�U��/t��>����Z��ɉ\NC��B�����}mHI.�R�9�G�/P�[�놳b��\d$�v�i�b��)n\��:��6��0�n��R.3�!�� ��hˀ(���ڇ��?Z~p�K�$J7���ms8��W�e0��>�&�$��@�໳9U�����NBB�Ң�Y�@�N�8=L�0읶�� {�m>@(�s�z�� ��P�$�L��|t]V����-�K,�Ł�gJ���`5�A+���IRP35�D����#N��H�)��6Y5aj1�h��&�6�������{�ˎ��aw\�*k�@2%�n�!�L�B�5�)i��S
�'�N���F!b~a.��L�������Q��]�X��?O�7�wA��+G<U�����]�]꠺HJ��n
�������E�Y&���y�q�((����p6;}�f�I��d�8N�py��.�c�>�҃�N��٭=��T%N7��^6�S��ﮮ	�r����1��b�Jx�tV�u[�L�N�YʔP�zf��{�Y�TP��z�M�I�0���m��W�udh���:r+I�L\�򿬩iOl�|[X����a���gw����ާ�����)8=�t��L�U<�\�}�����s+�	)��ٗrh����oq��+���n���*z�f�Ͽ��Ⱦ��BU�O�2[[1e�Y�j��)`Ù���r;ZH�ď����߰�ody�tz&=/��Ha]uD��D$P���o�T�Zw��)�>�_��tO�� �10�I)��V�y
��i�Uڈ�c����)�:N�^D��D��l�/�ζ�n�K�Aq�]Q�@*�/-L���c+�/##!4�����R�Xxza�}�A{9٬YS��UMܗ���Iq~�G�e$��P�c����?���̑	�	׃m7���@�	�,�5�9&�H�̌3ڙ+`$������ў�
�@$�a���Ƀ���Nm�k*w_?TLY�d��ɭ��^1=�J�%��:A��ϯ�V��!
�����h ��gD�^�Q�.�G �M��ꈋ��Ɲ���S0Ӓ�ȈO������6�R�!��]�'Mj���� �vך��D��VTWO=;���`?;'��S6F��'��G"4�R:��Tc�i&v��s��F�ߑ��!cMX��䨥�+|���Еx��#$�G1o:����s��0pA����_-/p��qJy{xC�
t���0��[���j7��C��s���E}�����7��܀�#��9��K��>�-��/1�]�:vc�h���,:�M!��o{V{R��#�%w���37�6iZ�0x�bB�G�\�WI��/�,D�vu�O�v��0ХG?[���*B(R�Gqg�C��)�mʙ�y�'���Ps���Ԓ�7$a.��TeG�]��ίAB{s�lw���].Q�/.X]B\�-�֏ad$����`��l5��n
O�J�Z^�5^#,������!"<��er�K��d����-���cE>�8�CV?U�
g�>\@QYۜ��K�L��ȻzO�&�g
$z�;v	̎H:4ا�#��m�gY	$bզ���̦r'N�]�?�C4q�s�dp�G�����D[b�dM���.���q��§��uCA,��y0�ݻB�/�2�Vo4M��ڞ�T��A���g�d�}֬��IZ?o�n:��X@���E��?��i�VJ����E��&��~yb]�Qz�56`ohJ�債��xy��Pu']���o�f[�[�ߙF@w�6��3)��Sz+M	q��L�:Ax����F��c�)a;(�686-#����Ą�r����Z�؄:f�͸#o]�r��Y`����h?�4x��u�ǧQ5Rw���^�s+`:�'������%,��Ɖ��د�
2g�\a��.�ʌ[PV���d�ē�ϻ����'��Q_�Bn)~7�>%GTܷr���7���VV�-0j�f/#\�}��4�)I�go�������Ɓ��e��\*W�=�����C�.J[��楌�Wrp�W�s\�3
;~��|	읕B���㍆o�܌�.��Vy1QP
�$%��Xe��U�_C!T�pF�Pi�~}+؏��t�ڭa�?s��o�T*�d�pλ�G���̷�����:�B%~����g\�7, -���=������b��n kn�xd�C��F�q^�M��	���V.D��1V�ɷ����\g0�`+<�7��*{��БN�{�2V�N�a!؊dC�Մ$K�.�>-�"�/qS�����R�%$��@c�����ݹ�߶�������Γ� g�d䱫F�4��m��%y�:��6hg���floxzW ��zA=�ό�Yn\udL���a�%R!��U8�:7t���nՃ�o���챎od��՜�-�~T7�	K�	�+��]��a���^��5�3)���;�3A��=t��֪c
̧޶�o���J3UI
����!3K�S�(�ܷ���/��[qdD���n����=i#Ab-��/�Q�y�R+�����9�f���{:q�-&�]f�M[ -z���	h ���G�X�⡦,P���3R�G$��B�T����:3�8.�Qf1_��=��޳Sn)yU-d���l q���4x���_G5���<�,��y�H2%���K�EH�Bk�����y(�.=<�J_xO���v�h�a
vwj� �V��pקih2�����[� <i���d�.��1����RѦ��;��Mq���<��l�"��V8N�m�?-�o�1�T糣k�Ʃ�aO�JE��ް?9�S�7��&ס��h����1 )��ϋ!�i�/���a.���$�#_�J�!��Bc��P��a���`*|�+�G�����#��@j�����p�l<h�򕊉�N
|���綠��n�v�����י��_y�sk6]j(U�U���"z�����tg���"�/���E��$X���z�c��Շ��w�t���-6?���.��䅥MZ���1a������aP���%��#�(�e?�}�b|�QfP�[�8j��Z#�-�J�v�"�24a����5��q� �S��23��0i3���6F@��� a��:�(7u��O��Ӎz��Z����֚r0m���/"rJ�VM	#��
(R�Np��d�8���+H��|�Ϡ�3��Ul`#�v�@�JS��H�ӏI�~j k�@p����+0�h���f�:�y"ۄ�p�gS���5���e��H#���SLn�B�8#N��wN�9&M���\�R1Ow:9�q�$�v={Gnmtڝn��t.�}酰�B��2f�54��;����=�n�XܦCt�C5�J6��3r�|Z�z���A�4����$�uϻN�
ؤ���a�ZT�/��X���W���E��m|�i��OCj4��L�D��K�\K��˥`�Bڿ�RZ��`�|����ᇡ�����b�Z�%E�e���PfM	��+_x������w�[I���r+�`�{�F�w-���H~�t�����w��h(��!t�H8]���W�YY=���92v�L�	;�X����&���<?s3���eC��!�.�|Ü)���(�ʝ��gw�8�F�x&�=�1h�r��jRM��l~�����[�b/��_L����K�l,%�SxE�7� 4�&k�!VEG�q�Ɂ�c6��ͷ�WY�)F�Wg��Z{GE�S�����W��hc�7-�!�m\h����YW������j�)�G.�E�[$����͋`Iy«fPҧc����"e�ܨ�׻j6�U��ƨ
�٘���o6�%#�e�2�t���ji?�  B�]���d𑕧����9m�M���n��#��2b`��Ԝ#�V�YM��{�[���Sj<W�'�:��W5�x���I�; �:���?�%㤸���)C��4���>��&�#>�y{Ҥ\O�t>�u|	�۩��w�(��{���u�f6岙_K 
���w>�'xZN�"ى��V���0݃���[�zAÞ�^4� 7�9n5�}���Y�|l<�9�<W��W��E�"ε%��߮��qz!���O���v���m��1���7s���.�G�٨�~?���N�J���NK����0��	4��Nv?��rE�qO'ͫ@:o�93�ڂ��!����r�&���d�dk��8)������j&K��r���O4D�Fx�x���Gi,:��I�B�t�JX�'h��5h�w�Mj�F�b
�͏ɱDl__U�2�on~rD;�x���m��M<$�],Ї;������#�9������UЍ,�KNy�$e�Hsܭn�Yy~)��c����B��3�_��X�Z�Y&u�=pˍ���,d;틌��䍖��>E:�oo��?	��^El�d��\0Eh�T1c���r?�'��Z6�#�`�H=3����K�k�`�<�'$FS�:�*�Zj��@�0@}]�����~�=��Hሣ�敏�L��B��A���X👴���W�2��[���oIi�Ɋ}#z����	����E�:����V�»\Arl:��H��˅�E���˧�;3����9˼�Z�˸E"������^kZ|�H�`�nn�b}T*��X�a.�[�Ǜ2�/u.�t�;(0�%��X����iuFs�T�@SVP2N�utz+&��8���J�ά��A,$�-�@A��G$S�ߕS�˭x��J{{�\!��!��7E�19�$��?V�)�7t)b�hJ�A�2.�_	ix��f��Q1�8'�>�^.��Z�LX߬�'���yVw�|ꐧK&x�0�M�{C��~�=o���H�!6Qy-�� MɶHwbU<��;&��I�z"��Q �Es�V�|�!�K�QSňRq�Ex�#��;s51#�b���X#`Rc�2F�|�PPA���q����a �lfR��QT��ت��\�ȃ�ds���k�V��iƦBs`��.����W�)�btZF��2�}���yϑ������� P�����46�L���&���mգ�3���͚1������*��N|����f��I`@�3���#>��fs$�_/�Ы�&�r�����C����/��3ؕÛ�z��a��-	&K�GK��xǢi�Z,sw�����'������	3� z�{�ʋ��t8�� �`���/x�� �J�3)��K���:Abo�8��
��ti��_|A��b�� ��u�����/}#�-��F�"�����ٶ�$abH�x[��Ù�"{�D�2���h��������0<�=�6�Q�)w�����F4��I�C��$g_��$߈��Au�;1ܑo����$!�E��rӣ��^9�6�x����d�RF����7k=�[�nD���5��+��^�y0�# =�-�7%a�	Op�bO��]f�i��V��A�
�$���T�Ӧ��k�d��h	�#��v�w��P�\8H��|g�%��Pk�	"��ZQ�Rep�н�0F_���U��`-+^�2�����	%i'���n:��.��WD���"�0c�8����0ِ^��x�N����s��`�pB ���&=�	@�����ª a�����h���nؿ�/d�%�4k�a���FhR����/T�a*�~����$��؂K�����7J��k	lg�o��לG����F>Z�e��F���!%ʕ"!��x7SB,Zt�������N/"G�Y+��)�_��6���h�����iNsꛑ&f3Ԍ,�h��0
�������:c"ѱ��Ԑ��h O"n�wݗ���;g�yٔ�˼٦���5ZQ�qZ!A�C4WX8���J�e��]�{PD�tH�~��m�D����gg�n�$�l�ŅX�5�u:~�
m��2���y����ﮑ<Y���������[Z�Ԗ����v�c��qmم:��͡����D��vf�s�-1[��*?�8mʫ	l�BU���U��7c���5z�v�;���CǠ��V���@�����I��G�a��	�0_�z ���x]]5�B��p�i#�V ���%Q��a-B\/�~[gY�=s���΂������Hc*���g�y�Y�� ��z��}�V ��1r���ccs�Xo�����߽�wǔ�N>�W6pz��S�Tњ�s��Cx�� ���3=��	�Dvb�3f�����yp��d9�oTq[��M��Cʺ�$2��j(�˂���m���!6�����P�*�i����sQ�"��9�3��]1�K"��RSC)n�����Ъ�����"*Xc�`�qhǿ;93&��TR�P^���=Q��T�0;���N��!�8���i�<��(�*5cKw�ƒHL���M���r0������[�h�[/^Y�/�ܾ�a�W�*��ҩTdw�)��}xM���i�̢'ȳ]_Qf1�g3QV��T�"Lg�y�b|
�O}�S�;b�|X �맭5Ç�e-F�>���=��%�*j�ߵ��"Rk��a�"c��h*!�&��f��}��O&��1c*y3r����*���йE�g��N_�kS�7&ģ�@�5Z%)M��&�:�\�Q�o��|?�Ʒc�1;Ш[|���g�Ū��T� �r����gUkT�Ҁ_L¾9�����cJa�N}H�Ϲx'R�m,��/V�Hm8��l`�Dl�yɈ��W4�qo=j���%y<C����mQp}>���s��S������m4�����%�h����Rv�&~�C����R��ܾ� ��監+��QY��[�U
yp�ê�Qw���& �u���)c&�j��h�cnbo���	��M�5hQ�: �� ����<&��w���%k�(@t� #��-1��(��N#J:m��Y��x��#�������i�w�Y�x�����Q'��x�H��ZD��f ��T��	>(�e������=IX��_^�����=my���������n��V�9��r�O_��"����׮z�9�҆�wٟS��_ II	L�Sp��ﵓ$�%�D�����F�؞u�`��.=�8�&�$���d�n�z��w���Dz�S���Y1�_5|����a�T{`[��E
 �������G\�^�]�g�i-�����j�}Sg)gj��1��l���̡B�^ќ�~���8�7�
�B��\��wY�ǜM�Y�U�h��X��P���	<��|�w{<����B����4%��_۶����ݼ���X���ƣ縅r"?�=�QX��:�i�Z��œ.A�n��:�R���lUD3s(��ɨ��=�e[�CQ�q#����R-e���Ƴ{u
��:����-��t>[��[��d-*� "��N]��e�a!���6���57��Q��cwC���Y��uw�5�G����o
s������>�T����H���h7� 01gM��T�ɍ�
D��'����_�cY;�=.*}%E��j����"z��ن�6���8����fX2vwj�T�-9Wշx���93 ��9����]��<j%q+�P���Tw�!k����S.ċ�;���|t�i_m�y@�20cNU$b�r��H��e�O�1�JM����&ZN���󱂍t��GA�S�<�.��?����@�9�F��J�n[���I=G��eq�l����c}6���L��������,mVfА��:�C�/�:�kȼ2v�(|���hA����_��(�!�%�����V����V��[��-�U%	ԫ�����(�*��^�l���
�j0UF)����K�$7�'���R�&-��������'�"��z2�o��Mfҳ��
�Vh�VC�׳-���lhα܍ʼ���	Q�T�CQ����Y��� Vu�68k��1�f���1cn?@�nL�[�g+o)`\�����0��*�[�R]T�b�jT��j�L��߄� 	���՞��G�-Cڅn5��"A�Ϸ����H�u �M!�?�(������(���d��̊�A`��L� j27�m�ʮ:�2l�^���<��77Ɏ�[�~_��ӹ�Nמ��>�RH��I�oGj&>Gv1�j�G��� v�)�ytҴ�Щ0�MhVT\I���@��Dݡ��}RÁ������s/Ҕ�����^�\m�*-T���
O61e8-=�fF�+Vi��f!2�n������6�5�WKe�I�Nf��#�E�K�-�ti�H��Yp-�N<���Z�-l�u�$l����_"�u�~L�%�{�q��UaN(.a���į��7g�ɇ��,CY�V+���bҏ\i�c9�(���F_����%$�0���n�>�&���{V`�,p�/X��;&�������]��@���<qŵ��Жh�d��"'f�T���W��%��D?����F_��XZ� �)��%\�ݵ(B���X�U�t���~��͖�P�I�[��b�G�@���,���Y�"r�#��l}��9�@����q#]�!���(��%���3Y�����1Rz㘂���V��
t�5�:9��=�)r�Y��[�Ѐ�����k�N����[������º��<�H�g���*��$2;�}h�5�{��)Ŗ��T^fa���X#�,M_6���';�Gʉ��S��l�Pz�;�������A��{�3�A3]L����CjF����l{�*�����y��~d.?yʮ�[�rŢ���֬ɻ7��l���iP�'���s�����Go��gզ*pWL9̆�-�"�~K�8��*�yO���;�ا��Q���к(���o��Ae�>��
�iH}���
?{�k�y��S<=��)"Kn����S�l®e�Xh�7��V�o�2����!ߛ��v+�L����؟�>2�U�,�5�fCl#�G�28����Ӟ�I�̓!c4��c-8�[�z�����.�� CC�:K���aX�� �~)�Xd�c?���;8tk5J����:{Ӑ��aM��	e���刿�ǡ���17:r����*�,�xZn��D������"7'C���@�Z�z���>�_.h��)�Bq�ȼ��kw�/��(l^��p���]2�f�ѷl �����
�Xb�3�U�8�M y�76jtn��@�b�C�ұ~k��`�(f+�QDgP�q���)sT�0�������9��ķ�g
\|U�� v8"n�1�:c4G�U��w���!��7K��w��ۍǪ�E�v��Ҩ��Z�{;��dMͤ�w�~�^?�)"x`�.O=T��~�k�U���;4�MF��t�P/��њ�h�([�VDn���M�{�A�uu�=g���[H�.!߈d4���H�l��\R���Kӹ�v~E�7iBr�-z-�*u ��Лx��]���p���g�wa��Iiڈ�ߗ{������9ü�)n�{��=�$@7��C���� o��|�ۙM e#�d�`v�NdJ���UQ���ÿ�g�q��NZ/'|gB�@�#�ZX\�j��>��beվi���=�rT�[��U���i�Y����|3��PR򖖶,�y
jX9�p���A@ ̹�<�Yſ�Q�e���hq+`LE��X���w)���
�^�G���I2#Q3	zT�ۛT1��{��_�%�V׺D.u-���>�P�t���m�)�(lo4)�݁��wWƣ$���v����n�~5aE^"�ſ��)Dh�
AL�cw�'ר�!&s/�["E�VV��:�bo2aZ�*���6����z��+�&]�絘��8�t�S�#ߍ+<kE���;���5l~Y���؞Ub�׈�7��� �9C�̿p6�x\T~�̸���Q�d`���m��+5�eX]�u2�Î�_���7�U�-��5����Zɷ�g>+a�4�'lB{�K�l���h:)�/�f��ŭ��Io�+7edY����b�zk�v:�W0�8o..�أ�R�B�7�Br�ݥځD<��<Ƽ3�i�@I��X�W�q�n��x�A��ʜ�=�(=�j��g�f'�Fn�TT���=1��V�EZ���v�I�N�0�6��cr^4�yOY|I�{b
�Fo����b
o�)�w��@���E�` �V�����C��Z�5k��i��V?�j�#��bJ"P�SA�0�X89GCh�##��wԦ��G�la�7og՚��SKF��s&یu�¥��P棖��L��nD��a���Caq�B���3qʸ�-�v	m^!	�]A���6a��7<~�ՓcH`[�D��O\}Ӎ�P�H�T�y�:!#a�:g`�ߐw����3I $a�����ʉ{����Gđ	4E�Y-I*�0��-�0oO�|����|�
�(z��J���d��,)�̼�b��s�1e���v���wSe�(sJ�9�e�dN/�#�ޝI��4�������L]-��O5�5��#R��������uٖ�Yݜc�����X�� Hrt@��cr����J6/|�,��b�37�<L��6�F���� �)�ϗ��&�<
`�>N��V�]`�I)��`�|N�}\��jq��e`i��|�>]�+�`��
�֤*p5�m��g׵�6uv�n�)*\� Nh]����U��vo�� ��hs����0��r�d@��b�
\����' NՒ�"���l#}n)�><��&�i�$��oW��B|�w�p�u�c��Y�(�Bb�c��l�P�0v��NN��qm/.fS�:^�d�H7aȷ�O"���A4��:P�;��Ro9E�u��}X#�����L:9���.��%L�?t�Zi�����h/l�E��?2�< m5�X/ֵSQ���ӓ%k� �Y��U�f%ؘ>c���4W�c:���Ɇ��ӽ
�x�n��~�3,6�X��L(ƩZ+���A�6Ut��/J�"� �M$���i�����tͷM��	��f�l�$i7q�!&"�2:9;�Aʷc"�1�(%�����Ɵn��L��<�TCoS:MU_j�ua�G͔ܯH=z4g�{6��C鳐A7�4τg9�C�$Bt��2�ޫS��l``0�L��Eӄ(��r07�������3p�f��TX�̢c�I��>a�.�4P��5LɏU���75.4qO12�����$B��P҈vy��2ʼ�]�s�%�56^ t�{�l?��y�� ,��� zب�W)����1�>��_3�t�Є�?����v�)��bYI���u���T<L�I�vso�Zn�Qp�_�cP��5���dk2��	}�.�,&�XwNbǷaV����Qа�y�?"�r����csI@�b�x��_A���&[^�Ѳy�����ad�:�����MA�!k���F�_W]š�������œ��R�H$���/����b0"�wɒ�񽛡�B-X���C�qZҍ���e��j 5<+�l��ߊ+$ �����ٴ�0l�g���M�V�����!��Bq;��:��˽]�Cw�5�l���!��KM���P�8%���nj6�/PO��k���2�螎96�kc�e�^ڂ�q��k�ƥ�D/��r�e
��[2�t��1;�#)�ܧ(��sX|�cwo`��cA�Z�[�9l���#z�l�vxR>Uк���Y?��>Ƣ�o)qR-{l��n:�/2�z��:E���K*!�*�\[��9�TQ����o�P�+_͠�zm���zPw#Y�$����QP�Q�B�=�0�:����2�h�n���Z~:1x��>�r!t��' �t)o|܀�y�TG<��QNy�y��x���f�<ߎ����ZX��V��jNVy�����33�|�G�����*��&_ɃN�#\`��E�|�T��~���"A�K�A47���V�/����J�x�Z��TVr��]L�!�8+À$�����R�J��Jb+�U�4���ɋ�^�R�?Cw3���G�T�:�ZQ��A�^��VGe��ʇs$h�7��`��,��ĸz��ix��%�1���i� ��og�9�ߊw�:6�2���34��@Ɏ�ܨ�:���7��×������0W	=T J����W4X�L�^�5S���	q�v%*��?q�="Ϥz�=��=����P���kX�T�B9ܾ�8)�'+N6�Zb�J�2yd�R��+9�~�Ƌ)������%��=a[�3�tR��#AN�_kE�_|<�:��J��4~��O�3�x�ߐ�3�d1�ȼ4 )^���d�J��Мf|�{@�j��j�=��DZ���t/�,+�v�\���D��f\��>p�c����z(�n�[�⇔���\�`����y�}���cL�P��<"*.�o2�8n����O��P�q���9�|��_�ص4)r�MT��`��X�@���qL2kʀB9��\�p�?�����B���z���Ԓ1�Ƽ��@6*ʩZHaI�r���tȢ,�=�a)	t� Si	D���<���kFV�/@G�7v�����4�`O�8H����L���c���>��)�wU��,b��'�F�׶�|��
Â�(�����	%P���ۖr)� ���A ��幂���@�d�}@�U�7��vJ��q�w�I�Gn ���XI��D���$I�WT���&��O$���%q4v[��Lr�}�3V�ݏ�j�hSԋ0��ɁSn)J=ϻ�x�:^�{����T�w"�.�o����A�j'�b���8
g�el�~=�`��B����>m���X5 ���z��z�<�`}v,��O���M�~��;��#���%l�̡9[)E&�Q���[��r`�`�����W�;�#����1M����qʓ�IZxa���S�:/ ,�2ym�������x�+���{��01;��)���T���e���>�~^W��М��XC�O�0��p���'��x��N�G��tn�&b;qiX��3C& g��P.�A�b-�<�{�Q��]e盨��F{���rV��v M~6��,����d���ik�ݩd����
.�<����޳�X\�όJ=l�~W�\I\h����Iz�v�ФV׷f��"��#�V_��� 96s�)Y��W�q��V� `,��&���#�[�z��}�ס�ϓ1��R^����t��r�2}���������
����Y�HP�Hb*�<s�,�~���������!���Y}AP��8"_Z���2���q5�.��N5v�ֈ߻� �|1A,���Y��:�,�O�jNp�4N� �.�Ղ ��8D��y��ՍO:{�w�̶9�DR�n q������`���=P�Vؘ	"��&�#�u���>D����@JƗ(�A���=�� ���J���� ���h�;7r��K��"�}Q�C)�H�$��%���ry+C���8LS�Ũ�ȡ�|טF�o��V�N�ਔ����)=B榼����])DY�6���<���T;�
^���r���R}j(R��@N;����@���WsBZ�.��S�sb���%E�ճ���H n2�����_<�N�2�g��%쵣��eQ&��A�$�#�u�x1<s����C���+��Z�G���� �p n��F3q�~��p==$����gμ��@�h͋w�|؂��<���@�8G"DI��-e7��R�ȭ6��so���7�ѿ:Y��=2�Oo)�/����I�<8<�o\���m��g�5!qIy�a2P���5�?0r���iU��F�B��t�n�K���_���s�Z�~�%�5&s����?R�Q�VJ��1���aJ7��˅Xl�fy�	�L^�ݹ>�T*R?Կ���h6|.�b�q��v���-t���x)��l��4U�e v�)ʫ�J���o
nZ���V|��E��ɢ�2�6�g<$���)�]	:m,4���6�U���"7*b8@a�\�&LY�.�5T����x�YM� �wU���A�n����#�B�Zbz�jS���0��Cyc�J�t��/�����H��,@���X]?$?
L��#���y��T��sI���ͤ��iMxJ.�x��T	��n�fɹOY%{r��A�5X]�S�Ձ��8_����WO<i'�>�t�%R�,��=�V��\;L�b�/����I?{a$!��	Q��8����%8��}CյS��1	\�r�CTJ{�N���VF�:"��k;�
���"��R콇�M�ݻ�p5�Y$}��:E���3������Fs-�eG#�ؖ�N�#�?���k��֭"��r��Me1#���AC�p���2�K7`�m�(��MQ-N�	z1R���aׇ^���_�C������ ޷^�i8%�<�jDP�X��ޥ�����<h�-�j4���?����1�O#��gQ;z)����(�#;��m��	�POV/�mr�ݯ|=L�dÿ��8���n3༓�б�xh+ׇ�+�5R4`:_��.�}P'D��e
��>J[�A��{U%����B�~8�#�˃GCd}�b��_.��e��)���|x�Yvz�c��X5���ߢWy�C+��?
�� �yY���y�zT�����Z���:�xN��&���跗�m���F�1��N+$h�r@GH��s��R>�4<���U�o�#��i�ǰ����iߛ�څ�|�]�����|�*�qfy����&�e�Qmr���[c����M~㘎z��+��Xo�|
���� ֋��S3��ۺ�Ek�Y������TL0z��'����|�L���1}��)Nf��pq��i�6���zdI�	�34�V��y@������F�^��Z�[��i��>���|�3p%�Y�I��I�ݗǻB�g�y����!.U���q���</Y�z�a���s£�)��f(�z�r��ɰ�����Qy��F�k&p	e@x]a��C���rI�gSK�.E��E�ϑ��|vc8�i��t%��q��>\�8������`���Y�^,�������^@�\dmWU��}<���V� �Dy�s�N���{F��P�g_��Oɇ�⁂8�ѫ	�Z8����r��W%�$+%�q�;��<	̴���Y�o��"�O�5̛%�c��"�o$���j�t�W]e#��(�;aA�i�
o����O����*Ur���3O�O���Cg�Z�qʃr�ͻ��V3_����0�d��Y�y�d:62`5,~��S���x�Wz�d����v�@�5�Ӊ�+����GYځ����UH}LT�n�2e���`1@��o"K���.n�з���P2a�T>l���2��|8������iZ���c����^-��t��s���|�F6^�Om�;�8]��Z���q*���d${�k���%�hd%Bp-Sn����z�L���a\n'����k`K��#�{7,۞��~����wӜ�����l\D0��"�s"�4�ݤ���G��*�{%�n�h*E�!Dn�sqČN���SqL*�f=�@ԋ�*�"�Φ��B�q��x���&O��X��Z[��I4��|�:�9=ƿ�����| ���/ �}'فd;�D�9�Ho���ENe0�r���W!�Ԫ]sN#�������MPZH �>6AZ~��h�S��O_`��s�_D<��iZ�	�W�`K�.u��.�/W��#�\����e��'n�i�R�j2� /�� ����� �@�Fn]��I��l�	T�S�1��3��_�3��s2!Ŀ����J��+[�� k�sC�.�NJ%�r)�s�^޶52�,�����>U--��U���I4<=��HK<���RH�.��8��K�����������Iٗ��^ݸ��F�ţ^%�̯іLȗs��������F�pA�k�k4�ks�φH�����WO���$�i"T��j �/��#%o�s���e�E���2^@�� �{|i��ӫrܳ��A����yTL�0���k�H�n�|L�,q���ޙ߃	��j7���'�:L�(�s	�p�#���\qX���x�����'��	�Ө��@�^R9}���ةB�p:�<�S�`:�*�����b��t6�sN*#���Bx�Cþ�W��p^*��6࠙���o��xeδ����t���u��$0}���H��� pf�z7vx�"�j�&^
��.���*�^����'��o����a���R@�yiz���lí�����N�Gt~Iۆf�@M�9򖾧@�o; ��X��	(��[E$���uD� gCC��-���d_�yN[�I�;dv�W~ع�/_��0׊�<��=�;�b�o�P�q�S#��@Ǿ�+��br�M�_����Cz5�,�1�������MX���~�����h�׮/��R%��
���:ood����Q��g�ތ��7�
s�4du����_`��z	SL�p�g�]��7����#7��Ì�v��Wy����-V�b��>V\�psx���X>�N��(r��S�ˤR�k�+���}| >k"փ�?��0q�����5���Z��DŒ���vWG�����^�9my ��m�/*y�$�\�Cew���/A1i�Y��gυ���6�+:���n��-�_R�;����Z��[UxHRK)Z�F���r�(a�aqX���˵�*�o��~���h���@�NC�"<����T[F��ZN	����Y`A����S[��3��,��h����٫}��^ R{Q|;�ޡ
�����dƂ�����WO)�ʂ0~p,�m� &�}��HR���������|�l�`3/��3*�gP�-�G��M��?\4�>��uz���+T���"��=��[0}�X��Ch���#��>�V1����D,�S8�����L;��!��<��k�&#7��~�Y�:���k��d����D�����)�ɝ��)(�L� �:�H��B;L'�X�y�3��oB�8��K��x�̣!,���5�Aj�.7=)Xr5{�y�u��W�h`u�=^%��G���⭟o�we��3LQs~$�0!�BFDS�#%#_�&�D�>L#���ӫt�'�����A�y�فV}ə�B�6�������0�N�*���a8)���,�x�Bzܽ���7�w�GE��<����*���sF-�z6���In?�M\�#'�o�E7([��*���5���7��u1�m��̴��z�W����zGAc�Y�(�}�a��\z ���i8�`��O9j�#�yF���H��3�6��9F�R>B���2#��h�#�}&��׉{��M�+P��8
�hZ��bk)}	�)���c�'X(�a](����r���h�T�*�!�M��>��U��mA[YR�B-.�j�^�O;���V��AA��Ns�	T�qa��+�z6�a1�� �I\v�YϦ,�y1u��l�$���h���(�Ea+.F=H2`�u���:��o:�~>�T뼂*n�oh	�JI�̩Zh��d�9fU�S'��v>D��`�S�E�ZAK�1�D���!5pm�pYfy;��fx<5P��]B ����J���s��y�L�ϴ0��hN?�܆h�&+T�D���[�Lb��p��n�n�9C<�
7�V�J�������lC��6~3����A��t��s���5�>��+6K��� �)��*��TY��R�OI�}_N���Bo��������w�`�ƿ%���.����U8L'b��D2*O�I��ׅ�*�!�"uwo}�_��~�m���\��h�q�Y�~:�&������UR���W"zZK��=g�Y����*���$�h�ʍ/�o1��S�T� m8��lJ���#� �9�ڏO+:�h^@��dSș��?���!ii?x9|�c*6ak���Pzog,d�X����]�Z]20t�KC�J��9_���t�іMA%�AW�֭�_��C��Պ�Z��!(R��3_��qӟ,�aRq�|%�S��+`�$-�z�z����]ࢰ8)%B�f6A٢��ls}�V<�ZVF��lo1vKB�gaP2�	Y鹕ޠi0�bb�N1�{bڍL��q���Ʃ���Øwx% ��ۈsK�Q��߂���2����ހ;�W����_�	���������l�����b'�s[W^��jF�=�)+jH��1�q��$��΢�Z7-�UE��[|P�yc����8@!���aÎ��U�*�\��}�{�	U;�U��rf[ٺ��r�h���J��o4�ӈ�ޔ�[�k�)��X�LCZ�S�L�o^^�	�װoq���*�<�0�v��5���j�Ɏ����xWю�t����d�y�$y�XLeFg����dB�G.S?�C%v����FGӖqD6��{vN���� Ր��MNOb�+Eh����*bk�|��?�&b��9���<��p-�Qz����"$ro,�;��+T`��'�����2�og=�w�|����폈����dO*�`XK�~���h���"�Rz��x:�\�D07���⶗��b�:s
����/J����_�����un;�;p! ����B�%�/��6B��"���{RX1��4� �S�sHPn���#��ה��c?bH�٥���UM</�5���43���\(��g�{��Ȧ�;���8�w��p@}fG���-+����9��@�GO�fHڙi���V��#��'�m�������<8���`'k�3�ʅ�w���ʼ${ ��M<���?6���K�Rk��
dɃ�h�s\b1���ܙc� ���Bc�e_`�G�)ƫ�fUq�FJ�+��K?�G�W�o&4 cI����J�7ơdB�i� jP�QY��)���ت�B�V���i��_�L��:�L	�z��k���2��H9g�fC`#.E)�!=2���x����U���AL:=���,���B���_n�|н3��
MR)����3�Lp���:F��w�$2m�-��x�D˟|�_��7U����#�!�MK��(]b
�?�q�Va×n��D�#�/��zbon V�У��>s���=pW.%���N�nYt�T!����_J������ZVE���#1s���D�Y>k�W9E2�h('Dn���������\�S�R���4ߚ���\+���� ��k�:%Y�*����9T�Z	��������GY;bO�>c�W�R�L_�h�R�կ�<��l3���	���+��hR�k�R�� SH��1u*!�e���ɨ�O�QkE �\�=N�1P�=��>Go�]p�מ�-�r�2�0u(j�3���"�_�I����%����'�Q��%wF�������dM�J�4�a�Ē���)����w�Tr	\� א����spvG�������a��|�<Â�!d�N�!���o_��?tUE����'k.3��茘|�T8m��eH�=��l��A�:�'{ЗW��NT�@2��\;�s�Ks��r�}��=ӞC�m�{�����J'�=���� �[J�q}��K�d�׫y;[�����|7�K������t��a�"��f�V�<1�B/Z� ve2��)��p@�?)����.f�"ڷ�Gzz��5���9�<��rd*_(�����;#d��1����X�;�Nv�bf��
�Z_jž���A*��$?����w&F-ؘ��]��0n�Lϧ �γ����+� ���N�}RPZB�P�����Β�K�KϿ㘰虓�_T�*i��d�	r0�U/'n��+���̕�tp��|g�D��5�4�%WD�b�����$a�?uS��Mer����/��/�a5������;ik58�;�v"�/mխS2��Dr�uP)�iɅԱ���[�_p�ǰ��yb���M���.bO�XƉ�Q��@~Wn�w�'�S]��=����8PNKJ��Xcwy�4"�]�Mȕ�`� �@��:���^-a`'I���GcX�c�\�E@��X��~��4�m0�)���,]����;u�q�u��� �	���F�7<�;�6�]�V��������xy�r�!��E��w�o��0�A�JAX����]��7vK��]M�G�j�[�1z�/}2��7��5^�:�gq�ߞ/�����_h%���6���wc#����,I/6��9+�����&���^s[�y��;I	��^YS)��6vAu�(t�� ��&C:�h��D������B�EZS�8��}��솀hhhW��8a�х犚�n�ڤ �Ə�m6��i�g�,UD ��溍� /����������7L��f��nӵ<;�B2H��(��Оz&�yPܻ��b���U���Ⱦ�;NX����d�m��{a(U�#���0�fe�q�0��^z�V�f��K��gEVpt(D�P�x`'�&���*4���ɵ=�y�Z��4Drw���]�HG
���j�/`.5�}
����P��]w����Bl��T ��(0��l#�#��E�[E��
�)o��C��]�O��0'���i���:&2�+�!�\���\����@���ɲTz�����/Ջ��Q�z��f�	�r`�I�7��ȶ�,|���;γx�6�T�M�2���vV�n���{�E�C��c�������nn)�*Tq<�?�@3~�8���1�N�969\�*�)s�!C�F
sU=Ķ�B�k���HL���2�~��\,B��X��;�	>��f�2��^��(f�b1����X��Q���˩T��
`Y����6�d��zD/��b��M�_���d,Bз8z-���Ͻ�[N.�J$m�#���}\���	:��2m?G*\WE�'�M��HV<D�z���u�_�Ǣ���[<�b{q{���R�#E��T����Q$�_-�@��h�wc�%O��^ 7HǺ���Ȕh+%�>��<�f=̤0��J��ڀ��j&�V��w��іrl"&P��
L9�{���F1��,�?Ñ�)�~M�
��������,"��3G��R���SߩWDv��z}U݀���p�wE�d�!�mี��)O�f���	a�cv��l*?/;ӿ)���W�@�nI���b�*��/a����c��Pn���]��~�> %�Z�9�#�;���)`��J���t-i��;Pl��%��."��?�����^���^1��2ꌽm�X����7�=�z�~�8�VD���G�m+�L������8~&�&ei��üЈ���K	bg��=�E�Ez��T�v������i�x)rD{��`F>J
����L���XWod��X�a�t����Aݪ6��;$=�/.�h_�t�92W��>����#H����ԅ�=J,c%	a&>n����aJs�·7��I�gMq��!��ţ�1DC�����G%���B�΂Z���7�96��Y9Tp{�7#S��7��s.gqkVwFL���}�Į�x�>9M�ĕ0�����8RŘ݈�vy�UP}U gR7���I-�e������LEN����UrY��W�o��՘ǽ@��sp���˙��D�g��/���e�<Ho�ـ����M���Äx�l�+!��!�aV�E%p)�JV�g�ޙf7�ѷR_=�S�Jr}�����P[e}��4�Ѻy��t��b#���=փ���|̎I��)�j�S��]�y�t��{�f�v�5Blbj�!Zp���1I֐+��8 �p�������gy�+����,6�;��l����{�Ke� 㒟fa�>�r�XOz+5�J� ����GQ��R��D�2�?�cR<O����u����o�m)va�5���Jh��%�R�0�E|��tA̛M!�|ׁ�'���nPc����Ѝ7������m��;����]P��`"v��y{bQ�\�Ia�e>��b)ע�
i�&���!��IGEU;�s7����`�*���\�*3���7���ı�·��xV�ށ�Tg����75e����FF7��x��g�n����a���Ɠ���k�K"lz��_γ��*��iJ0&�21�w��"�!�*vQ��1�@D�@��y�k�t�߁6����O�#�1
v��#l	��� ����d�zT)���v�x��\������F�-&�3�3z��"��n��^�s�V)�~ ;��� M��[��Ub�������Oǰ�
�~]hYU��yl�����qFxg����iD�?��\�1��r��iEZ�SI�\ݞ�~�	���Ր�+*4����A]��p�xX_��YY�{aO\��88��9��#�N�G� �/��U�Mջ!V�EE�)ߌ�b��Ǿ��b��5[�ʿ
�Լ�s��E�_����UT�j��r��5��N�km�����U n�����Z:��j`ҭ�of�̪O%�S��S�l�,���n4�tN�H����EOQ�4�<�SR�JF@�����Β9�6��2���d$-8��P̳�W�H�_b5,����@�F�H�����c09��v�
N�^�����9U2j�qv���e�*�%��	�D@,A�D����E㔴����Лz@YQMb�����ޅ��#�)�Κ�񗘈e�iB��AF<�qcl& [�0�G/�n@�dI�E&��� }�u'g�����ov�L3\���U`E�N�C��O����/�y��:4����vl`J)���Ԏ3��GAA�?�����r?%\n�n�0V��n��4����o%�]lBg�˫?�f*ўt��bDv���K}8rƪ�h+�W�+�8��~�������!��< !$��]a�}�r��>#v섰hҐg��D}\X����E�U(��mΛ:%�%�k����4E�ю�6Q��'j�ɋʹv@l����`"��,���sĘ�y�pG;}I>�T�rQ�'�%�҆��n�������s
�Z ��@��A�QA�j�2��"wô2����Y\m����:z 
���pWM$ޅ�&L4��T������ɞ�LZ^�f�*Y�u g�?(�E�Q��4U8�"�:��d��z���g�߻XλN�9�$�J9^��aI�el�j[��}���+�C+� ֋z_���;����o<@ק�:O�JJ��6���g;��J����\�
�D*�cH�}�	ֽ���COq9�;�BA��%�×X��� ����+���wSB�5՝���瑚�__�?CYs�Ϲ�(
d(FϏ����cD��:$�IRv�(�ӿU��eQ��bĺ��Rʻ��7[�+B2P;��pAR�s��[�H�³m���|���U3��B��#��t�#�硉��ųte��je.��;�>��I@o��X����ւM���a�����b8Bl�ſ�܆�)���M��.v���P�a�P��Q�r�/rY���L�}y3#����(e:����>v�w�M�����X|����m�`w	����.Sz�-���Y����ӭ����֑���W��u��z/D�-��2>�hڅt��q�����T ���xdN�KE�u����TP^�q�Ȫ>�_�d��-�e�U}�dX����]�#�M�+�Ɍ����o�I`@�{s��y֧p&=/��H&i}.�L6����T��x�������C�|�{'L�cZ �����$�x��[�u����;5o��N�b	0�jGQ���6s�����s�ڻ>� ���:2�Ter%+wA��������笳:��_�!��%�ه�]��Ù$f����7��Hz�[P�m��p�s��N�J.���]�q��e�N�N��[pU�P���2�@=���*r�W���B� �)u��¨�b��|��|!�����-h��j�޴̥i�t��@ xkS"r,1�@Qcm{������H��<���%�Gq�ߨ���%����a�\H����R���m�3��f=xtuB�/�-(�F7�P}���Vv(�Z�,�7gQ)�7�䓪L�:�����v��@� L+�j���m�+��=k\�Y��:��M̠Wph:I ��U1��;|���a�+1+ft���� �+�*c\N� �N8Y�"e��NO�R��n 7D!�����~V�3�-յ�>ؗ�x7'n>f8Ҏ��B��MY�J2�aI`O�y����ޤ�����&U;�ʉ��1�4�*�2�S�՚p9�%�t(���<N"�:O;��e��l	H�ȓ�i~/&d�s����DĀU@���8���о�����ԏ!�*��+�dg��Lp�z/��?��Z��w���GP�lS}�waT���&�,��_2x�8C_�o�D���s��=eAt�����ˎGB������2Kf���̒�ZQ�� f��Sy�4]f����� ��h2����D�G7��n��ђ�<`E��������Rc"^��ub�G<r���[{��BX��Nn��#q%�^ߪKP`�c��
��R�T���=�>H0�:���1�w^˂R��v��"�fP=w���Cq(��hT��������E�]�����@%[9�Jl�q�6uSbS\޸��X<^�Rw��i�`!su�X�/X�[��T_����́��x��Ci����J��K��w�7��y
�ߞ�s*�#��2��&����,v�����=RG���� ���e��D��)�nd�o(,���^�
�E/����{�'n�߁x���\��Y�s5��#˳���+����<�_\";��g|m�~�"H.��@����hb����5��fm4��%3s�C�4��B�y���<�!Iqc�ߝ��5?ӝ'!ɂ,4`X��;]���q���ۑ�P�S��p���%{�>_Y�=�ޢB;��@K}�"�S�w��U^�Ea���w~����'ofi����`uB!'F 	z����5"��\X� +j�J*��Y�#�+dE�*�n�ŵ5K���o��k"EX�7���*f���[���po&N�Ư&����E�dVVƌ 3:����ʄ48�7�U��6��������` p��۳��L�o�@�7m%�GX�=(ݸ���	�ԁ�J6,t��妽'ۙluz!Ss��Ҷ$g�C�}|�f�ܕ�Q9B���Ϯ
���me��X���,�����1�g��?r�eF$���^蓖F�6�3�g�'�7@1�g6�9�U��N����6O�����!�"��'b2��Lh:������~&�� �i�o��b��k��sk�����&�����ck���9�[���G7ַ�PfFt y���CxA��ʶY�N���?��^��2iv(ਬ��%{,x�	%"ȟuX"�	3�Fk���:~�����H��1V"*�̹�w|�D��Ѕ��hdM@B�!o0�� ��3�#��q|������~�T��9h���Y�ʦ�����L�-dmQ�-{���N���u�x�0õ�Pt�+�LQ'.#������ѫ�N�7:��RDהN�2�5[t�uƄ��;�MmM�%B،������(v����ۏjp��YC+{uA٣��QX�ߜ�1��~v}[�:���-a��UZ�@S'ig����U�m����:g�Hg}��c�<�lu�;�ZP�B \֢0��$���Yb՝.E䳮���d�����1O�d⣗/�>����rP^�}���, �����w�$Ki��mUH}����hgQ��$l)���]��4��	���|�žE��ӕ�	�m��I�ێ�e������C�WMzj2��5�{�(>�i���<�`X����͓4�-q����	g�k�>؅����ש���ϐY�6Q�m�>�!��E�����������5l�5b��)�rƏɆ�dN����gTz���y?�H���n�6���"���t|�.q��肐�9h �)@��օ�ٸI�Vx*��"�w�i49��teM\�v}���3w��|'m�VI��/k.l4S(i+:,lϡh*����$�G��4�߃w}�Ԩ�H:�L��уTӲ����b��V���Krr۞K�t�HJx�,�LW3Iz�c��R�1�&	� �����`G /1K�f��4l�b�6l��v�{���xZO�Y�	h�6�k�U~�:o[@KJkZ�0 �l/R����4�����`�'���	|�L1���Xn�`0$�"�-��x�{I�0�Jt�(�H�Pz�]��<<���B6����#i�NO�\=�81(~���������k� GkJki�y/�7<��kD�]�+-�ｵC5�J��ӄ�-����N��{!��@�)O�P�2ޛ��#U2"�I��Jo�v�N|Fln�l����2�~֞m@ ���U��3h��.�[h�|����F�:�B�l�<<gm4�z!��<�T#`[ԉ�	�J6�|ۏ�����	����=\KwF)��p����~�g�L[�*�� �N�Y{�ǥU��VC�:��О�����[����ҙ�0���0@�Dc+�����M����|ဍ&0MVU 6�-G�I4ȗз��K��Cɖ��S$���K�p�`4c�}l�\����&qQ0�������qVN˯h�;t-����V���ߨfI<�$9���*N�`>��P�'���<&������$ݼ�~l��j�N'�Wgu�^%30	���&G��Xn���**$�ޯd]�L'k��&�7��4yȷ������7�>����l�������!�ڗ�5YB�(�?�i��O���?�j�	,-!l�5���S}�
�n�nG1�_y:3\�
�1Ƚ7Q���9����ݦYv7�q�{�$�%.(�Cd�ˠ�U\����ŵ1��EN_��>�S������M� ���X������^$�`K�x�
)l�ec�������S�(�����\�E%�t�eI��Jpl��'��^XaO�m%��٘��$��E�~e1"'{�ca%l2�^��Fq�4h ҃��_�s/��i�`q�KFD���Z��aީ��T�n���޴ݽ�+R7-�D*'f�]d�j���< ��̟�@�M�`-<�~��>���2x2��1(2mN�&&�� ��SnB�6����'9�|2����`��BB�=L�cN5;;ؖ�1��S�Q�ڟ�9��l�m2Ϧ�~Ds �l�J��7Y1��B٣x�#�_ӏ��?6����X����;��]R��Bv��ݲ�+�r�;2���2{��~� ��n� ����z#|˩��[��FVs��2x�i9��a�Q��Y/��d��G$8�,@��N[&���אZ��6�UEfUƆ�vk�����ȓ�P���BUxE@�U�d%x��ĸ-z7hY��y���ؠ'�馟B5\xA���ȩ�K��:\��k��+8?���+v���VQ�\D|^є����(.��# ��qu{T��-v��7!���' 8�MW�&K6�&� i�B˽[�4�B����a@CG�_��WH�ϔ�Md�q��~�A����}�a��~���Y�ywJp;����tp(iVN�yr����bS-�� 7*��SY��+T������}+�,�񩿢ٛMcV�z�����2��>�F�.�\@��ؗ�HJ���忂G�5; <lt7&w`,�y4c�~H����|�Ͽ�Ee=m���{W~� ��u�,,�7l�"�2\���% !I�7/�TI���p"�5����Hl�gW��}D�_<�ɠ���ͲKF ڶ�uz�N�!������y��F�Rc�.�fDT�4����b�?���[0;|N} ?Pn���f������dA�u�u�]O�+�tiF�.KЇ�����$�ĬP�cWl��qê�>B��;������3�g��Q�y:M&����J�?��t����F]�.����pt�~F6��-?�Е���+v$N�LߔF�*s�F������]b��0���f���O|�o�M����
_J@�B-��>�]4Rj�ƾܔ	5$jN4s�������F2�I�fZ������#l%��CT�(���/�(M&�W�?���"����#�a��p%b��Ч�����=�J���5�s�#��yR��͕��:Q\3�� �o��(�S�ǒ��؈��)��D[5�����0�$�f�����AHji�g4qq�=�.�s%F�Ӿ	��/+Z�������(�1}��PT�ق��L�'��q�~�y(�F�7մyR ��O�����`ʼ��̥�u�<P{��a(y{O�8���@���0��eo)BcG�Q��vs%��
��P-,D�y:jߧ�7��"����~�0���0Z�-����Y��x�YW{��6��k��W���^��d� $�i��t�Z��G�e#0nVc�3F�>¿����of�D�m) �}�z�]S��Le8H�h�mT\	���n�h�u���%*��i�	��3p+6��qA�+���ʖh�J�3x���z2͞��/G|��x�����O!����
Fx�cA�_HU�	7v�������0j�#��������B�H��r�Z�r��⭝����'���g%�el���O�Q��-9�Љ��i^��愷�&?+�`^�_��DYIxK����}�Ί��,�^]��_Ƽ!��dP1�Y�ƙ�d0��n(��\ϰGg�����O&���qF��Š���ֵQ^B�>��`���)���^:Nhr8�-�d�P�S,�(_k�X�R��,G�<W��o�U�δ!��M�]�b�ȷ�8�t
����Q�!�"P�Y%�Vq^8K*���ğ���dQ�C��Jw�&oP�1�܍��U2�O����a������M����0( ��T�`umn;��ASL����R�j�#�bo�T�(�z.�(HR���Y��p�K�*�7�$����4n�]�;����KRvUe"y::��_۲u��@���8��n_z���XKy:)�B��,�8��I�kp&�z�/CЈ���윭X*�r��܂@m#^������E�5'ƥQE���3��z�3;���O��6%��ŹF����`M�b۽b�E�E��>�bMB�ם�<}c�S�"��f;D�@�Tk���/0t��530�����2%#'���;���> 0�f��q53��?���dA��+����n���ӂ$"�IX=o��5<)jmq�CBt�L�z)eT�>� [U淜���	��@0�N~w����͓rzk��'ۤZ*3��F���<�#+u��c�Q��A�"���i��.a��L�Ẑ��)��o�ރ�B��t�ᲸfnQ�d*�}������/��j� ���g}���4�\���C`��e�ڋ�4[eE�W#­Q�`���X�]�/�T� rʒ��/䭓8�\gy�=�Ź#�K/�9�.vLp��Kx�P61��3ҽl�8��ǽ*�´b�j���3�!�&y��χ	���
�JEotn��IX��C�?�e����`�:�R_䎄;#�%9ud���W�%�h!8�q��ynP�F�����\�����DK�q#+'�5��O�t����]�S�C��fT��
���*9�@�\:�\Uc�6���헣B��� �E���)1��ON6J Ũڭ�*rV��)��Ca`I����$�$���t^�bn�h&m�+���ԩR�@�@�J�{*��_VP�:�>uM��KY�g�|E��Ə�fݙ�m*�Ĵ!O�4���-b��g�'�����[h-��Ʃ�J��=��P�L#��\�j�$1C�ʍS�o2.�%��b�ӌ^�g?a��S�e���E��t�QN!vS�Fs�J��P6.��T
�ѹ}��B���?U���p�}����X��K�d6M�	�<�6"�G�5U|A�<n�������@��K�_b`y;tV$ݦ'��3�d�N���T�Զ�C�.t��͉K�e���6�|�Q���$�6%�J����/��bY�ժ��+aRߎ'������y_Vr!\��4���)�#@��*�EϏ�ds=/4)��� /X_�v�/���֙N��Ǆy�Ah�QK��#,BU��-X���aZ{_�M���Z��:���/"�߿)Vpq���,>���˂d��no,~HH}U����z^������g�:0K1JD�ı�O��}>�M����ȩ?�p6�UO\$%��|����2�j��J ������n�P ,�]L쟬�M5��,DzN�a	�`{T�:�[��
�{��z�;�n��
8�  �,Ɯ9�(�7 ���d=��Mņ���X��O����L� �D�4@�x����k흹F�\:>�ɽ�� �^q,Z�!f� �������"�g�����R�ۻ3�1��:�m�r��O8wݹ��[W@�pY2hP��{����<�3L_L:Q��'5bS�+(��a3��X.^ضSa9�6�䬃ʬ���%��E��CP���5+ía������*(Z)��4�F�Q:���h�g~��6o�P��K7Abj�5ğ2R�pWY=����~��-��-�L� ��TZ��M��P6�'������X���	���?�:w3=?ޫY]�Ls�B���3�t�b�.����l-7
�Vˢ�GMT꟭�3_nixn��PrHK)�6���� ����z�T�F��xe9Q�/�<�H�|�/��W�{I���ݑ�ϭ_�0��k�쨏_�TS�������f�v��>W�G�9����ǰm���z��F�?|��Z�ߐ�v)��9{J?�i����P�Su�k�~>ι��7ƴ1 i��03�����k�Dt�",��y �]z��q�����r���_�]Z�}M�
Cy��{�gB�4%1%I��>w�I�*�?jz|���dsG���A�B~��?իs�5�T�/�3�:��*G��;�Z�=��`�&�H����2>p�W�(��y���>[�e����1�@0a��=�]�|��TT�z��)���*b5~�D�9o�ϡ&�KO?�D3�˖�	"��\�ٹd�r}�*'��fv�kyՎ�ɾ��E���Z79�:�4�"4����H��`��&���<N�{�S2l�����"2�t���0"��yZ��ˢ}2h�������qH�#��}v�^��ޮ�!g�,u,�=�6Ax�:h�'�����%ǫ-G"��בuk���8Z�d/z5�Mw/H󇤊�|h~O��y�BA]�����w�Ӄ;}�0����r�ξ�x�s��c\��F�	�23��q1�r��};�T)��ߑUA���m���TK������a�;j�I�RE�
�V��䖂`f��
�<��i�����S�\5�\W�U�v�h�Db �&~�� J��H�������e���*�O���5�p��./�Tл���!.��fZhrv�r>�{^Ko���D�M���i/�Ԙt��d�z..�g�	
��gZg&"Q�b��O Cb�8��2U X){0h)�Ȫl����e��wcw���v#���槎\x��j����:�}�E��!:�u�X���X,:���QY�A�M��]a]u��3T�/A7�x
�<h�c;$�DKx��L%Y�����$`�j��f����8W:��g:�����3�`���O0��^윩��.���	FЄh'��	� hX(�5��4�����;�\��&�Y
���@	�G�MxvHל�2CV2���`?n�px!4#�p����LX/���灒3��-����h�0�u��:�����տl�aa�#2V�}�P9Qٍ@YĊ�@+G3rW���wo�Z( ����j[����`)8��S�}�j&�0)Ak*�[�9�����	���c)����S[fsq	��[�*�1B6U!�-.�T*<���}L�uN�9#��& ߐYK3� w�^b~�� �T�.6�'���F�ԡϱ@�M��q��[c�������Fq��=l����W��V9�  ��/���B�b��z�ο���7�Ņ�Ԋ�Q�ZWů�e/*�S��,y6����=x�<ά���7�<I3 0�2zp �6�L|��Ϋ�:a^J�Cwz�k�f�(�C�r��� V��N�0�qe]n�I�/j@@�Ug5P�(�o�/F�K&䲕��#20�O*Hoۤ- ��g�IP�O��W&��IZ��(HVk�<t�9�%[]ge2�FB�}�D¥&��R�UV�f/����8�&K|������ٯ�"�Q�sǟo�����6]�0)�f>�"���80����ɱe6��j�tT+���ӦxW��3_�� �C���
,�!W2}+�ڿ�×��>b�/�}�}WC��7��i�����6�p������E��>�a�u'��|�S�s�u+��Q���1'�,���F�5#oϖ��M�(clhn�xL�`�}>Mc���[���l?��D�me5s����T�J1$���s�+��j7��B�C�m~��>�^*�����_��BgD�&/��-��eT�X�/S�Qzh8���;f]o�\�EYE��}1�G �hh��łli())Ų[a-�7]2���ʘh@H]7s�U�?�[��.\8��Y�0�E$c�M�9��$N%6�ͬ�v��	�������{��o�jӲ;��O�rOcH���v�����UM��vC�[�!D�~I��$.'�x�i����On�<��ͼd��w�fN��k�2y����!0�*,w��~O$Zc\�H�#Q#~{ [.|[T����w	y�!�������+D�ey��4������[?�&f]V���r�uD<����w�`�h�R5�1�[�,a�V�7��(��?F@�.�o61���A�!� ���3 5,[&k#L���f����5��,f
Me׹�ϰ=�~n>���s��x5N�O�|MJ�+�+� �Ľ�@�W�'h^���RA����T�u�YM`�,�#�č�v0������R��T%�<��ܢ'A����y�Ʋ� ��~H���R�o���a ]��d�b���Hi�D����-��{ޘ����b�?�q�����������a/et]?ܬ	�8��a`�6� �Q�hTG�������%��5�[٥��P?3���"f+�~a;���j������pj�7Ӹ�il�pO^
(�ץ3�oB}�z
W��ƨwY`OE-v���Z�)�;���L�@�_�,��c��)����d��xu�]�!= �@E��'S9�;�u��s�ʒ�%��@�� ��Q�=U�\D�k��ͤ��o�O��cո%;C܂���d^����/��i��Zd޻AJ�r�|&j5.�f6�o��:�VB��߈8Ⱦ��v�����Y��	�{G\��9}_�-4y ����#<� W
MQ�!�(f��&9by���qc�f�iA���G�R(�*. ��[�Yƫ��qu[��S�x����������L�P���*6�l����G!(��	��{p��*��3^��j9k����^:V�c~�>NfV�rK�F����D�%�M$��ѢO{=�"���hyj?�sW���0εPdhU�S�������|���8&��l��`���9��j����%�]ԿN���g;���Q�@O�����A;��M���Vc2�ϭn��i~���$�+V��[L�kZp� {6�)����g�\/���$��Ŧ�Z��Y��cG7|��Q��?N�@�1�s@���P��:*:���O9k�ڠT�(���syq����U�s����d�}���
�|B����!���@d|p}VU)�ҏ���4���C.2��֮��~��R�*T�F�0��V4�C��(�̋����d�BH���y�a�M��Ӳ�a����O��{_�[�D�\f������v�`��B\��S3

nl�`	�̨Z���M]ӸI��P('Ն{J�>�|4��ﻤ��PӾdS3��P�nA�<+�` .$���FW��y��=��\��:���Z�6Uҏ����TXo�r7�X��P��B�pk�g���䶴�k��	�,- �4y�����5�' 	C��6�l�U���6��B�_�!����T��$�Ks@m��y��^]�+e�(7k����x��l�/�q�5���R�j0N�6*g:cWD$�ޑz�l%b[�bQ���*4�~rC;�{�!$ST�15f�i��x>k
i�!@����Қ��\���!E��vu���OO,Ʉ9H���>��n*���	D�g�ql���J=�g�q�����}p?����(1M����#{1�D��5,�ލ��7�%�{5S0�^���C��-��k7�֜AOX�z!I���|�q���|U��{�7��{�'9��M%[ɽ�X%=Kz7�!���j�!3�\�Rh��A6�Wn��-�熆z���R���n5�A�q���7r��+3P�3��W�&���Q�}�;���+HI��~9�V��k��"��7�I���N�p%�����]F�a�8��d�����F�)F�i윫��=2��׽߯�CfI��$ �[臐�s���j��X��o2;$/��X)u�Dnn3������D#��e|���؍Ғ�$:��3���D�㪴��
�t�+��J�1���c�@��4��ו.���i�A/���/ښl7[4�h�j�c�jw̅��iW1�K� "G�z�H|Ԣɓ��d��I,�f�6.��IB��υ�綝�	�c�
�^�I|�pNfn��Ot�0y��Ϸ��{\H0��p���d�M��+�p�ȩbS��eX�TA���~PN�U�d�@}��`���@�Fp�1�Қ��F���(`^ag���/n�"*+�>q�����Iψ,�oe����6��`5Y�&S�\�t�3`�E�z>-͂�_6|�>yg��vŒ��N��5/��t�k�}�娉.��Z��{`]��C���C�tp��^@��v��8��ɜ}�Wȓ!���h�")�h�H�|܅�?ZF$�|y�8� �c�l�(t���g)�;y���]L�p6]�jA���A��vc�\� ¬�f}�m
@i��`d�^��	�k�<��h����goB�2%���u$R?1t@���s<#o����d;$����$�9=g�-����hV�����@�����7�ƫ�X������vM�6�2��6|�<�ĳ��t�CJ�/ӤA˚���1|�~Hʍ�21=��������)��jh_e���Շ��Zqv� �R���|UK�t����a+p��Ƽ���t%��8��M�*s�Ľ9z�)�Fuo�)t4�U�sbEf�4\�
RlJ�ϗm�M���|qv���
L�l����ir7��q���6�i��+�B��u��Qe&��@l������_� @�ez���Y�U��m~�h��.l�����\�3f���V��Ӛ�|���d�Ipg�Ke��.L|%/�KЏϖIM��V��������Q6�<2R�Fo�E���ϵ������P]����3�d��P���v�w������}~��M��
��Ɣ�hj6l�(D������ro����[a�K	.8��^�<�#?p�C�G��OŸ�����)2`���vޖ��@b��3紀JG�	��* 	���e��:\ȳ@Q�a����F����}�E Be%�K��̐������y��-�b�#�1!�AF��b�12'�{w�>0�u���k���9��8|>���ٰÚߐ��G��) ���ݢȚb~:ѳ�U�����>q��I|Q��akz��x�+�
�cl��?.����.c���]�'� �q
X'-�|$h���q")\G���p7[ed�GJ�������n���FX���$� �����s�����;?�:y��D��';\�s�A���g�E9 �L<�8I�r,-ד�08g���8�j�0*�P���j�����O,!�5\׻2�w ��Q���\���)\�.4�^ f�Vm��u�t�F�(34��=I�v r@#�CͦY��D+!~�>r��*��� ��e�"�׻݇L�h0�D��*��3�/�1�:�sMظ�E43{�浟H���U�1.H�`9�BR����?�P[-O�\-9���C[�o-.
q�#�cI��
�9'я���ػ�*��Ȧ��
v!���
&h���B�C��
W��D�w�G'�Kd��`����;�M��66ua�!$KG:�h�L��9�F�z���2t��uQm=�]!c���N�kT�ȍ��Em��]!��t��K5�E2.d�x��C��t��Y���D�,q�Z��5�U'���{'��7U���=DM7��C/,�'8��1�1_@/��B�5n��S�/Gy����h��%.q1A����Έ���U���b�x/�^���w��Q��J5qE�BZSL�Mx	�O���p�5��k�
��O��Yy�a ����6C4Zu�7V�2idG�X�T/�����"A�m͚:��E�H���+l���>	����p��޴��.�����`�9����G�/!�ĕ��>�.�v;s�����3�*4�n0���I��˰ZL0��#�Ij=�aB�����+C�P"ͯ=��;m՜d �-��
>1�n��Em�V�T�Uv���}�AIf�#1B�LPy-WI��s�
�����eee^-B۞�4%5=��<��h��Â�s��{�>`V�JV���"'�Y�(>ΏE�N��Ka�T��ͣl�W����4��Z�ྺ��5�&�S?I#w\���~sC&�����&���|�Ϊ�xW0�㙗����Ŕ%���W+����=w�m4$�,V/���������&^6]BK&(h�͝�H����������6���I�8�e�[��4��]��C"[\�� P˟9:Rl;�-��8���Hۆ
��pP�K�ǐT~������}Yv�WymU��VQ2��P'ͬ��Z����`6�J�6�אN-ء"w�.���LB���������8�ߊz�d���D�h<�r���ou�Ql����)��O�.�+�Q���T����`((jNI1G�?l�f]�[w���5��N��a�GEpH3�M%�����0��� �������)�AS�F�*+i�}�z.�WNIA80�T�әFw!5�?(у���b�Ȥ��vg�Md<�y.�i�@�_1yC�R��	{|�p�Wx_�_T����t^��"`�\���\�IN��W���#��� EQ��<�g:��f	�^ċ�5#�����
j�w�mzT��S��_�ǌ켞��D����i�0.�9��z�[{~��2��я��)z�K�A�;�i�cȠ=(�'�q��}�����A�J`�%o�=`���T8��ȉr�:a�S��1����^����ߖ����w�TAM\`��g��υ�Q�'�@�~�h�$3q�W�����I���/ >���\� �	K�����tS-T�Q��O9	|@���f����)�X+�^�9o�,XI;}^EG�ÿu��A&
P��y��q(����
)��B[a& F�l�DD�PyJ����ʭR�h0k�GF�[�q4P�cvPb.!A�ѫ�?x�V"P��poZx�c�h��ڊ��U��*�%���xte�	�)$i˄�R����4�p'���h�5A����ߢ����0�%dDH�d�j��t��A��*�m������h��f��ܬ~|�B���8�awr�i0��3�*�-t�w͓y��R���wM'Ř#�0ol��F`oIIz+5w��R��*��Q�y���?:
QO��'��CT����]7?#�L�w2�r*c�gG�s�o?��F�}��o5����d����8��k'�e��*�I��l��c_S�Vj�4��j��5�Fc�%P� V��M)�w�J�I}�.a�ԾD{^d-�� �E����K<Z��y�	_��\&,�0�d˾�$�?����2�s���x��d哠����&�ikV"�e���Aw���'���)N_�H3�G`�90ƨN�VOSG���'�Q�"4u�d+����@���h �d����(Mݵ��L&R��_Kߏ�xC� 1�s{)r�:2�g�l�iU�V	`������W��؋����D&�����3t��t95��������IY��$�z��U��cV�mV���T)c�R�O	�*��(���xfA(A�(�B`�\l�~U��g�`��Sa3����п���7�6sI(S^�l/`Gr��z�dϣ�d�|6��ؿcYHΙ�3�JC9J|�0ڃRE#���}�|�.�f��ﱉ�ۘ�����o�o���y/�VL�v,�H�4t��!��H�*Fl��g�~����ql��a%�l~_?ɷ���;IO���4-(��]d�N��0�g�����v����&�Wׇ2�!q&�|���÷l��<uha�CT�W�f�~0ᗷ�PH�b�:����:��>ϣ��0��Z�&��7Ț�YY�wt\Fo ��W����)��4>\ ��L��nE0�M�� |�A��@�;��
{�M����$��𢜻_��W���2���Y�Nd_n���?����^�?�6��wj��.c�ԛ�
�X��
}Qװ	7=�4+�,�,�m	�Y��[N?�61��7�:P��A���槣��+vZ]�fF��ɫO������x>�k����%[���C	�_����eG0����e�ݳ8Os���ȿNJܠ6�������.��Z���8��T�ϜO�-=�1c�7k������q�xjr��;4����X�5eE5GA�V��#�&jh5ϼ��|���7RW� ����ޟda�oS���Na6���1OùY9�\
2ؿ	��-�I!�a������������U��Ӂ��9��n!�e~�9!�T7~�b�CT�%�b	�'m֧�7f�5�8�Ä| ����%�o:��|��N��������,c襅[��5��s�D��5�bRh_[��T��R�K	P�5��r����0�Wq�cO�d� ����@��C�5̳�6�yX"l���?5G	J�t����ɝ��c�*��tV�m���&Z�z�jWX��1�Kϭ���a�h�$1K��9���D��U�8N�ʜ�*3#ms�XҠ��h4�8�nl	��ȿ��LZ!��!�?sJ�1�0-p��zϻ��#z�򄶬g�f��I�[��e����I__"�'E(Tyu��[O��q�`:B3�J�i�bˀ�b��I�ۂ�C�/4��zM���}in/c��q"��~��
�,�a���X0��%U���ۿ�YǬ�J��5�O<Z��6��i��zCyD,��?�q��ڞoi�M�.!�G?ZV�IrW|����t��㑏e�v!#�/n��`��?O���zkj,[���X"���]�qq݈���Z�Hl�K���>"r��.շ�4�n|6��q�`ч�oS2�נB�~_/GY��PM?�b�eK��������R��XE���	�;�;�RXB�	�.�}iX	�oE��Z��
��;G1���KE��{D�?�K���'�m,�#eI<�y`����ӑ	'H�B�p�o�0���o2���J�r�`�Y���������2aiE�\��Dń�ߎp��w�.�Af���SQ����bꪩ�h��}�P#s�ͨ�l�L�j~|��g$U�����I�&(�I�G����R����{�и��=���{�g-�Dc<P�
��>����.��FE˂�z�
E؟��;��8׮,W��f\hi�*.�l��֧}LQC�o`���F���B��6+��.��󱀄k|\�s(bp�
�Yns�j<����ͽF�5�~��]���-��=�������]6���&	0"��}F�n�i}�'<� ��~��� 3��j���g��*X�u�v@Jq�O�8<����=��Ih.r+]��d��� �����M~d��,| �-�!��� ��A�Rz��;T�M~�K�0���î5h/ӿ\>L`�.���Ȁ��_yV��̌7l.u��i��M�ЈA�O�������߭�e��ΗRky4��{�W\DyD�P�\~�N����Ͻl������b�)��6bn��zi������r���L�o�eN������:�5�צ0?vj�W>��Ǳ
��'B��f�F�,��?����JCqD�hoV�1&�d}��39J��k=Nb�Q�1��+�%.|���d:���d6�Y*�����m�e�W��{Y��E虓�h��}���g�ô[�S�f�@����۵$����Ŕ�{k6f�ɧ�Ĥ%����S�;)jX��o�����`t#n��	�j��?t�6STKZz��s������;n���I�V�W|�nC�k�X�����eC첼z}?e��t&O�������}���b;F{a�Y���n0ٝ�!mss��M��p9Ԋ���P�Gl����Db<���mͰ\a`�J��";\���  �X�dT������#|��ʁ�?�+����tU�hY����ʭ������ȼZ��]P!���,���G�u��Ť���A�f~����P��L�����`u3�E5�e	cpR7b�9�$n�t������T߄�iws�Jp{�;����`�z��x�Ni�G���+l��ؑ4�}�t%.��s��&�Zw{�)��+H��5��YN�G#���LCLz O��7�/Ib��.iQ��F�\��w��-1�t*[��j�U ������Z�c,m1uCzr��-��-~$�ܖ��JWĴ�C��>�p��;�<l�o_E� tB0Y"%*!���� ���Ya�U������ٙ��ST%���������)��O�nA���㡞b�E4����
g8� ���P~W�.oӫ>'�Q-E�,H@�� pCF2��|L]�#L�x��~F�S�3�����ø.*��D9J��,���g1�+��9���?�M�ܠ/�qm���w������V��D������Z�9�P�e6_�`a31�eݍ�BB��Y�/<�r����㮟���'1)ۢ�E��cP	����8�>Z��0�d���#�H�+m�;�B����@� ~�!��Ø��f�׳����=6���MʼL*��'	��������ihU����A�@�u2<x�K��4�w�>	��b\���b�%Q�#��T��,5��ʶ�g	��!(�M],��b*#�\��f��)�!`��Z�D&¥�>A�-$��W�<�6\M��1��c1�`X�����E��	� '�RW�E9.��}��O�DR��JŖ�M�=u)�Tӫ$�|�?��@�q����^�,a�E%��gid�H�b��J�dȴ�d�Ӄ��]�K�'a���|{�w�J���������#�s�G@SO���M9��z��W�U���Sk���Y[ˢ�ߴ�J0�L����^/�!W�	L�W���-�&@C�\��ⴳb���"����اd�VЊV҃'�u���HQ���~�WީB����r�V���9$P�K�G�TJ����}���"�fcc6��9#�i�H����eUSX�1v}R�$z��cד1.@�)��C2��B�S�i�?;D�!]��8�mN�����z�%D�_���#��>	�81i���<C?Bc�����>^�����+�)���q�O�OjJxʄ$��$�0#�tV��cD�����f
ķ�}��E�9W	E�wg%�D�����G�	�O�k���4�����8��̗5�ʃᴖ	�����jm������;��"g�g�gI�0I�cgp� hU�,�����k	�%���>Vv�8<><E��f�/HN+~��/����Јe�]��u�飀RT1"�*��q��#�	���E]��hJ뻞jkiK�w�)eoډ�ߢ��5��?�n�y0Q���9J����ꌿ�/���!�@%a��-z;���v�o�\M�:
�B������1Ɨ֒��Ro���-��L����Z�S4�h e�������|4|�,T��9qEs��`�^�U��ش}�hS�|�Aj��x��97E��i�F���$Ƽ�0sl��2��č�б*�+��\��"���Z��9)�?��BQֿ����ʆG��nJ�#w`���wZΰ"�G� ���+VQUX����y�P��$������Og<
C��z�8�eQu�T��992�����	�D��Z�yӚ�S�8.8�7	a�t�
Mۓ��s��	M��^�=@����B:��V�/1���=oC5��q�w�E�u�A�`����gL2��S������bn� �J#:�+E-��2-Ʌk�R�j�� �A۝�S���`��u��U�S!��2xT�3İz��3�H�,g�p�+�/J�4�~i���l��X�~h�Ku��0�bZ�p��,��a!U[ENN�C�Z]�z�@Hx�V��j}��ś��ά�E���Q{�Չs^˽i���..��"�/�	;��-k$��o�ˑˤTA�F5w�k�������tFI��?���eH�/@�9�,��� wl�c��OU��G�@y��"�D�u�$��:_"����b��"A�j���y�g�����qß�/�Px�i�¨�^��eI-���	a��M�z����MA3j}�.[=�_
�����}��$��~e�I�v?�l�6�V+��YPI�.՘[�2��V�-����L>jZW�о�U����Ux2-�u&�9�#D���2M����/V�9��z�a��#0i��Ư�
X�^*-�^E�])��BVe���裂��f��P7̶?.���u�b�7͠wC)ڃ!}0�\1��Ey�_�_o@hGI6&_ȏ�ܗ�&C��d�!O�������$�:�T�����_�P	��	J��Ss���:�A�Ǜ��4� ����[�~��ABt���8_׳2R�ʨ�q �߂y]�F�h5��(^��;�o���ޗe����l\���$�L��=���Rv�(?!� �� �vWO�y���ߌrk��3�-��|�rA��P��泆�8�y�Ŷ�����%�`��
 <��=�59J�We�`ΦF��	T��{��5Y���@�~}tϙ�dT4�%�qVK���F��w����#��M�D�a2�Ê�()NA���C�]�4�W[5o�P��Z��8�k��l5i�kT�^	-����d|��Fѵt��[�~�a�8y��"D����Q)Z�(?�[F���0�J�}q����S[,�;R(a�r���'(�ﴅ}Ɉ��ǭiz�,�:Vy�l�C��>p/�/9&�k=~1��)��7ӈ�o�Jɥ��pfq�*��,�B�q)+�B�; H�BH�E�'3o]p}Z�9�� ��>����ܞ�h���B�#�=4!8��+�LgNB���)�񔼜�p)�]�#�� �bF1���h��:_��F�Q��oG�My�ࣉ�+d�qp8�x0��`6V�G��3�����
������:~˸��_TW�9�)�}��!Ԣ7-Ĺ�[O� #���H)� iV�_��V�I��T�e1t(x�l�H~n�t<@EH12J����T�����ώ^�
�K�b�K�V����
k��	�Q����
2(�X�0į����H�*]J���H�]�Ŭ��R▇o��v=[`�����ϡ���0�S��-.~F�')��'��6U�������ꮐ1�bC�KR�� ı%����!;M���}8��'fCO��X�(�y��zcR�aV!���Wm�l͹���z�η��v�],��{�*�F��j�' F�8�5`G��~Q�m��f��W��C�ΖU�������Ě�]���d��.�w����R��@�ob��{R0�]��*ϫ�@�1�I��T��������pk}�Tƕ5s��TK�)Q��=ٲ ��' �)y�~=��eZ�L ���Sr>Bȣ���i�H&�ج���ڑ�bT��n��%��@,�,d�!(W�9Q� ۨ
�R�u	�F�+m'�q��Lӓf�g��h֌`�S�r6a=���:�q������]Q� /�0pJ9!Z(�t���y��Z�.�o.����l6^�P�u��fYLa9�FE���}۞QZѯ��1��p��B.68)�_�/��c��V��/���Uan*����X\�0���ʁ�Ȁ:R�n4yYv�\���''f��.���r8�s2�Ҋ�;�{?sDC�囕N�p�(����h+�k�/ܾ��������P>�E�t�6����%d�!�;%2	';Ԯ/���Ӌ|�v�ʓ���u���%�@1@)��v���$�g�����OӜ'�n��G���Q�4��	��O����b���c\/+��_p���6��uNH�Ot+���<�M��>��{z)�p�:L�8SO;s����Z朗cˡ�^Z|۾ H�Ǩ�]�aGۻ�^2V�(n�*�X�}�Јv��=}
Y�Cj�e�78�Rb7��]���� � ��h7�}GXq�36�{�U�ch�7��������T4�J؉�{&4���E������x�ă��S@��ӗ�(VӶH��������ˡ�NbJ�\t(eR��D���D��6�7%6�����ӉFL��c_s8>"��i�*��L���Լ�vt�k�Γ�rX�?���X������D�*�Z�ׂ0a/1��G|�m
���m�˯��ϝ��}���iJp��]:�J����]9y�CZu�tVD��;0R�ޒ��=��Lt��+���c������j�R�K�݋�i�C�H���@��'*�=�Ǻ����G<�J��p�V�<�/DS~Wbg��Z�((�B�Z�Ċ�K�� <����3g`�ѩ��9au/��E�p�ԋ�^�hZj�Ֆ>�9�
��Ĉ�;�U>]灣"e�xt�bP
mv|�AE�K��o���ɋ��ӯ\��
�
�9at�v�py.�w�d4�q>���b���U�?ȕI4�����5��s,�C)ۜ09�f��Ų.8I�SMA�NC_�.�*^��y.�涕RuIkn��D����T�(���iY�@���j�g�46zmW��^>�&��#}��xW��n�9:!�T(>q���|��`�e7���� R��ɰ�{1��/�]�|䅡/}�~�y��l�΂���=/�JqF
����ex�v���1%�b1�#a���%��*��2��n��V���.��kP�z	3��p�7s��|(.���S_8���Aݒ����tl�e���:�$����k&���3>�yb� ՙa��Xh		Tvs��w��.�Vfר�g�]Qz�$^��k�%��>�&�eD%�L�τd�vr$ ��"QmōT�5�3�`�7E���)l�c]�W!�17BwB�e��M%2r<tw!�x���]�~�Bq��8�g�,u_�0������t��H��0����w��I�Լ�j.��5���G�����!qא����F���tF&�Z�l�(K�aFߊJco|��DN^ʙ[>L�w��
<8��n�0����A�k�>�T��	�j f�Fq�`2tL��Ia�5%�*"����=���)���V4�e�?X�B���8������ӛ_����ɘ\qO�R�H��Q�4�C�36/�w��� ��8���L�^�k�t��a�'�8#�й�w`n��gB�1U�ϴ��qskF��τ��9�4�?�C�%?É�KS���.�Z��W0Cq��7��C���"��mI|A�h�Pm��~���:��h�ӡ4g�xu�ǉ�籵K�y^#|$�h_���
�r�� �g�}�����l��M&�����x�p �->F�2T`-;��k*5f�ds�}!J�.hǣ`�)w��Y�����&۬LL�le^-��YTrE,4���U������]c�M`x�ȃ�ՅᯊB߁77k�_ʆ�����'���9��d�h�D���ƫ#t]��n5�\.�����Sl�S8l�j1f���+<ʺm3��9�>�Y��1 �ةp{M�/��kՇ٩:R34U��ۊ�L�|�����+[�b&_�8�T���~[M��w�����/Z�9ױq�,�+o"�#QV���Xe���`�eMT��e���)��7x���X-�	��Q�,Y����(���c �,vc��S��E?�d��i[�ޯ��wV> ��䁎�`Fg,/63M�aM��r$��n*q���tU$�1n� [�r�Ʒ�ew�#d�YL>K?� �nä�ڔ)DR��K���bۿ[<<۳)	���H�kl椘!^�fN�����**�v'`�<Zn?yEW1�!̝]��
K�I.a+) ����>�¶��*n�2�C.iC�1P�����)�"�$̚�^��!/��1�ď@rr0��1�S�������O�5�^����uv��|ǖ�Q��K�	^���P0W�C8C�OK��djN���
�}j�����x5�"�c9����=ؐ��L]}a�%�de\�"v�/���@C����b�w]+J����*^����9��*���@L�\�P��	�Oq�a�	�Yټ�A�ۃ��Jx�Ol��e�RvcIY�a�R�>�9^ɷᲹor��L��W*��"���uƃ;���}�R:��͋����O ����$,�X�U�MI��r��J
���\��+B\��$ܤy���c���ʬ)���l�f:$h�6�8T��5���#��11��-vw�.z��X�seY�&�CuI��3�����Y�ᩤ���S�d���Pk�ϞS�a�A�����b�H�ܛ �O��1�@�v直m.�]{y��z�e�H�5���U�k��ZΧw��U�E���;��I�u�Z�
'��о�J�|9_)J|�s��ԃ5g��=B�\�)/���o�Ŋ�Kú(Ah�OL`��n���el�pA.bqN���Y^:k���0/"�u&G�;A�HSkn>X���t��j�l���I����=�6�Wt�B[��/(�ܤ0� �b����t~��vmSwhuQ����y����鍯�r�!g��{�=2�9*b��˂\sa�Z��27b������ݣ�F�0[D񟓾��V�eUUGab����"S>M��/5�'����s��c��H)q6�d��	S�
�J�<}�$�K��C`�� �����!�4���q��.�Ǚ@L�Bm0�	�o"���7��d���P���a5P���qlF��J���hΘ�kg}�>B��o���r�I�)�:&���m���t<U�IGB������Z�e��5��n�ޮjr��Z���St��k�����8�[�d�ן�CN�&NDt8#��
�-2�x��n��/s|��_n�K��g�S�U=��`-?L�6�k~Ɩ����G�&���% ���9'��ǐ-�;}*򅉁�iOQ�]���i��Z"t�5c��U��Г��a��[c?f�;���uy���ay�{Ǜn?���ڪ�����Ca���Xw?2}��FB+�!�K}�|�l�����;6�I����p��>,��K�f�����*�W�&��E=���}�ڭ-�S0��-l�M�@��f'�=YRֿ�>���h+X��c`6P��U����a<� �W�$4��(b�+zⴜ�����2	�.��erLս��]�z�G[��i"Mm1���C�I<A�jhD'�m���*r�2���ll�s�˧H��{'�4$���Ol�o�X۞�7*ޟ
�|���ON�������`Q�8�-Ƞ�d`Xf���&�28�q�c���WK�)E�Y]@ w�>85����\�� ��8%�����K���z�)��H?Y���}r�\���sήl�u�0�ҵ�hIobWb�c�KoZ���j���D����X���.��_ _��,[?t�����m�K�+�{S$���#M����~��h�"�֮xe��*��w���î�����pG���.֘ 5
�Q��G~�ң���Oq�Ke��ݷ��<�6sI�,T��d�<���@�����p��{��%~�s@5�j�	��ص�9��`�mBWT�+�ő��@�f�f�Z��o� ���O��Yx�}�$�t��5�z���p���=�/�=�)����p0uS�B�*
Y%W.��-��B�/����h�Fm�940 \�� ����]o�o��t,��I%5N�Ӫ� d���38���)i0�I�i�9�*^*'տ4M�zΛ�ڜ��Z���f��G6X��*#���U��cD��(ʆ�L�;w�?� Fc��7tr�>�jѨi�C���8�6X,~x�tD��l��;�4[w�D�$��<�&��OvI#�TmF��� i��ٍ@���4����1�72�vub��"[��9c�8�0�W��9]�d;�LOs鹥nq-vT�(��(:!R�[����>��j����X�m]��[�t�y��q(հe?�<[?�*���l[�|�g�L��~߄n�HT -��l�nTAu�Z�������B��p�"Pף�Oc�m_+�|r��)fQE�'m�쓅*W��eUD6;A�B�:���[�np�]A���Rw?W{Y�.���Wye�b�oU�x��gx���"�\?��>�n��ix�L�$����P!׀{�>�M#�[ �.X��c�/�$�G�6���腙�WWh��[aHKx�t�_� �R�N�w  m��u4�}�������C%�琻��w4�P�]�͑vh<����� �#��	���B��~_�۟q�>L$�žO�kkO��[(��M߷���љsa� �]�TbF��:�a�mv��N��B�ͺ �7��r�7�ԑr:,�l�q�R��[sw'�8&r��z��'ȩK�~gL���������	q�h0jb�Z�$G���|b+♟�Mr3m�lCN���l��DL�ܟ?�h�R�A�Ͼ�M��YF����#�漍f	��)ĝ��+~pi�(&K�M�y���D��Q ������X�Z�3N��-E�D�p�)�����Er��MaCc�@�.v��E���V(��3^��<H���+**��E��X���Hc>��y���.dS�C++���E���:�iZqTܖB���i�
�j����թ ��j����;�ˋ�È�0qA.���Ś�M���J&����K��� ��SY5�"��3�z�F�3}?�?�&�S��ρ�휎�y�Cw�Ԁ�#�|���%�<K)�{F��GN�]A2D)���� �]���V4���-w����O�k:��6�+l�Np\�����b���R�Dv&��W�L0>� q٩Rb���$݈���+���+���U�Lb<Б~����d�I!��O�`ԝa\�^Nb�Ӱ��Yqst�xp�<6�ćɃt`c��I��5m�m����l]3h�f�</�`��Q���Q�(Wp�:�iZ�<�<Jw!:V��rݻƌl*H
�w�j�������s��(ʡ8"��6[
�|pd��v@!�5D*lQ|�L�-�� ��g�~�S�Q1����Z�iX���� 3��a����s,�DԊ��xSm��z��̆N�[�e>��K�U*������/hsj�z�є�[�s�RN���pF��죘X�l������SB������&��2�R��D���9�zd�Z�oGJ�}d���6x�N|rc+��N�I�V���H�)���3�s"�"��<M�A"xOlkWJ����~��~'7{�ײ�9 �Nf���Y���������Zjm�5� 5��7�r����x�α��A;�x�5�h>�UAPg�8�(�R��#�m��o�ؕGU)�:^����/�礮����N����`�m�~~S�L�vg\����륶�Y�~)4�e����[�8�l��Zۋ7�ؑ����=U���%�#��(��0ں`�-�.���ض�Cm# ��&HC���J_�A�����m+ѭc�{z�)�̹n��v^o�[�̚��u����a��(�E<��C�/��8�O<%U�������ly�o�z�z<�3�c�#"mF�U��_KH��1��bbWmA���_���r�e�n��U���Vʺ6����i,���cʪ��*�ÚQg_�l	]�W����:l�dJqXR��AS�&�,o@�EL_����f�.��f�s��Mv9��aZ(�8�������hE��,�զZ3z���r-<蹠�y`��<��6�>(��Щe=�|O�����#�V`��]y贿�a�<��
�<��R��ѐ���Vi��fd�7SQFz�{i���n�牂_�Dp]"��"E��1Id�i�p��PI�$2��#�9z�h?IL�W���<���)���ߍf�h�9o�(K������&��0�6�y�QP��ĉK�J4�q��]��֋$#"/���0|d^;|�-xw�� ���4��9��,�X!�qt��-�ί�5�Qv��ఛZ]���2�k�&��fLM�M/:pa��ȣwq�����_R�"I(������7O��O���V����lF�b�Uj��,$3
m���$��.��_�,�����iBΫ��c}�yR!Mb`�c	����`,�����@ku�−<���դ��&���}|Y�+� ~�d)��W1��*λ}j�=��`oL;��Cu�l���CE�oerV��+�"S)��'�Dt4���9�8�8�t�t�W}Ԅ;�1&r{��;[w	�v�Y{0����LF�2^�X��CQ�BRswN����J9�"��0�%���0?^Wl�_�bR;��bA��r'o��E�Yw�y�����e�⽩�٘`&�ZC��~1U��?�����&&|�-H����t�����cE*�AM]�31>8V���G��!,�Y�x� r���M��>�
q���Y���9S����S��"�!;ۮL��I�~�0=�Irl��G����f�"��\������3���f�M�ߏ�pܝcD@���a�	�Ԋ;o?��x�"��%\`@�1��h���W��E}8^L��7;p�Rp�42ݡrz�C+ޜ-3X�w�C�,h�u���� �6x�m7->��YlYT4R���F����N�b��X{3�8��͙�8�~z�I��
��}�x$�֤�f8F����REo�B�T�c{��	c��fҶHH�֧Ŕq�t���V��:��%d@�9���!�g"����}��x%#L�z+��E��O�GҖ��bo�Fr3,72՚���y�����RͰ4��p�k�\��� R�a�>��]:��[�e ���mœ�s��¿_�P����Ǖ*lq�u�|ݰ'Af�m����{g�;�	Ҝ�4�X�K#J�_y�\�3]�
:�pW�s�A9tT+��A�e�ɪ�e�z��$��������{#�Fq��p��s��>�<iM���@�C���3!��H��)9�8�~	��ꂊs�6S�e��$�Auԁb��q��� �=ŝV�`=#�^?����'�p���b��@�~e�ɴV>�G�6�'#�FN��$.?�;������{�O�."�<�h��_a��B�#��1Q���n�D� ��;�V�Z�`��ŕ3 C��z��=j�_�K�ގ�tZ�3x���Z�#��vK9x."ρ�K��SB�b܁sN߈��[��j*��F�WkZ��X4�#�>�j۰�ŀT?��+Ex��9�VM?��lL�w��x?�5@�~e���K�%������*1m[���F�%B��m�]�vhQ�ȋs�k6��S�qzo���y�y���$�WI���6��~�2��w9Z�^��Ѣ9Ƌ�,���#��2 �@b*3�p!�.Lg�'/�#f�x�ڋ��s���~,�#*X������Lty�o�ܒ�|�r����y�l�po��ݣ�����f�����p�c�)μ3����� ��Ϻ�a�����5�3�W��Q�1���N�� :��'T5 ����#�����G�����M��	�C��v�ӟ���gu�x$z7E;��ȉ4���q8����3}�w��z����G�.E�I�d�׾��௱��@�Ł2�?�To��6&�#���%���;}��N�ie�
�+ďw�w
��׳5h��ah��tHG�>LS_;_E��Tؽ����⁥�gq��@�u�Ja�A�x�cZ
��s�ӶaW���\w�T*1"��e�}������U�Eh(CFޙ`��{ѕ��xQʡ�t�D/Kju���};��9q�͵�XE�����v3U>��;X�Q�l��r�����|$��U������Yao��7T Ct�lIL y�1Ie(�Ihy,v�&� ��WM��)�XDLo��M�oz�	�a�M�o4�q0�K�<�I�L�[�t�G-��#}ɯ
�>s�n�nk'�v�p$jǳ+�a���vc�eF�$\Q?jݟ����O� '��M�r`�s3H��U�b؉�G�!�j����K��3�:����W��<�̿y��t�L�_�f��t8�&��v�`��6p�����-ߍRfVR��[���8�Y��`��6_[^Ҋx�;������v�'L�y��󕚻�ծ�k���r��>�FϘ_(����	���%��?��k�C%�x���)���r���~hG3��z�9�:�g=#�൥�a�n�:�}Ow8�&
"�x b���B�#~��*ڭ�W�|���R��Mn>ص��� v$���a��˲��>ؔ�Q9����p��"SP9�]�؍'���&�"~
�^����/EO=���J��]L8�u7~���&s�K�i���Y�O�oǑ������9��@h����������qG�=���o[���
)e}���h2e�h�{7j�n.��}H�)o�H���t��8'z�5��>�(�e9���'&����r3d��-�3Q ���]�0��Zi+5b5/�;�l��!x�>�E�0�C�L�#�l�	]KTL�Ɛ�u#jv�*�u��#����	J�<4��qr���5V`���3+�B�&���y��-eD#�
����y���OO|w��S��-��G����IݔSL�j�z���S�#��^�w����^�p�a��~��UJmh�o�裵�A�(%�bW^�R-�۽�zh��;V���In5�v	��"��j���Go:.Ȧ�*ɔؑq7���jZ� ��-=-�D��y5
�9q�]� Y�`�0B���@��R�0�3�p]����6�X��5"���
���Q��X�H-@���F$�N��Rm�a
��[�8/H|px5͡������(����K��p�~���:��O?!�]�1sCI�L�O��*�Z)�Y����%�	�ȹ�q�}E�����*~<
VW��ɇ�fl{Ibi�9����hW
Cշ|����˾�V������K�^���7G��8�]8~4��/g�giI�\�Q��7�,2��r!�̟J���@z� �h����t4��y�+}�J�N-ˣQ�JL�{��ׂ���q���7
����ˁ�O������e0�<oՕ��m����Ҏ�줛0��f�[ș� ]���u5���Q�3��/}�,I_�S�,`���ݖ���7����r�4���̌d%�ox6��V$��]���1}�l-n�7� ϧ>ܽ��/p��|ta�G��-��Uq�L	j�I�FF�1q��`W����e���x	o���sR��Pr� S����������m��3�4����OvGj4WW@~앦
]�r�{'s�z��N(��u�Y�oʽ}��zӲq�	�L'�ｱ?��*[y1E݃n,K�,�5z�l���,@c�� ���	�h1��[����EK�&�+���Ñ��#4�$?}otX�ڛI^��\�VJ��������Y�t����/�j�$GT7�u4�*���[�"%>�W��7?�2����&�[{1�F����|<S�U2:�QFo��qp�VD�C\��p�%���鲌��E�!p�_zE��CT&0��S4$�0nɶ�S!i.��	�o��b��Y�Q�/�o�_2����"J��G��Й���/�eAϝ>՗�����>SB���b9C��Y��!��bH�¥��ϵDǬ�>��/���,*� d;����E��M��6<�k��aw�?�%���Z��R��I�kI�	c���J��@�q�PL��~(���5U�YV��	���ڦ��v�~�W��{�!�7XJ9*�+�����K�L'Tˊ��Lx����'�rw���hO�B���|?\�W������-��+�#�m�!WC�gw����p�����nnbN/i�T���	.F�V�}Yw�U6zk~DM,j�eȁ�6?�7�]���/ UK��a�C��U��-N7������Ym��=���r�'�-�ܱph^m��Jz���C�E����t{K��*f�2l��BJ��U׵��_��]X���9�G���Ɣʪ�:t'k�6���y���� ـ�XdQrf)�t)_��8�6%h�sx���wM5�!W3��q2�[�E���MD:ʏE�"�3��g7�7��%�C���^^�vz!R���Ie�v���	��qePmP�t�Y��m��\��vo$�����bzkĵ� �� w'Z1�=VV�cȖ~^(��@2�����9�(�ʀ�j��º��^�
��I����(?MN��+[�g�߄�K��=)�`̵_m �C�,(��<P�m@���`��T��^Eyʘ~F�Xs�=s�S�d]���oye�2�_n�b��6��)�,w�Fְ���ǰ�dUmU)Δ|�'k?��d\FA�ݨ�w����!���`�u�^�
*{���Ǖ!;�7���������A*nj��qQ�*U3hf���[�U�K���ഏ�J��oI�����1�QF��*N�$ߞf��.�.�l�܄�ZA����d������3jM��e=������Ԡ�+��RQ��a�#mZ��]��i �-��p(������� =���G����U��$�Al�v"B�%:��JD�hTC����:Y���ދI����=�WF�����@X�W���ja�ȟ��a���$���A/��Aо�׷����=Oo׾mR�A:�x�A��k-��%
�y,�_� u�|�O_вl�p(?;|۫5���օSd^�t�t��Μ�p��I�jU�Q����c��a�92�d^��)�9_���ɶ���2�w �+m������Vu���&��y��[X���roH<��m ����Jxz�PW��Z�N7E�r7��5$P�D��+z���V�U�ب��&,���$ޤc�#s�y���e0֔��K�LG�B�4�ﾯ�+"N�g���Kȵ�:�u2V3*�*��ڧ�v.*:0��N��I�s�+�d���+�B�򀋤��)	i��TZ��u[�i]x�e0�qE��1i�PI��,� ��r\vݜ~�p+(��_�����K4���ы��Tg�B<z!oz�0P��d~�q��f�M'�����lWi:bޜ1��ľ�+3Y��8
��i34[�Ŗ��y�c����)�0�4Շݜ�m6�[��l���C�w]1Ϛ^���a�Ɛ�.�'�6tÅY���\	#9Z1���@\VIpJ���!~�z�P�ē�]~c4}Pp+1�2�r%�JZ@�Z
 �k���O����NR:���k��+3�Ip	�-��rF&��L�)Gr��2��"�7�<l��$����6N��Q��q��k҃>7�k~�?�\w�:>��	��7�J��Ab�|Nj���i�-�p����p�a�D.�k(��q^h���t���vp~u�- ����)�����'b�c�z��"�ŗ�I?�����k��$����j)
d��r6���إq�|�H��JN�d2�;� �OZP��0M���u�}�T�$�#�	םУ���,ߊ]��}�G�z�ZZ7����f��l��d�߳��z�q�3M>"o����#v�7:��k��`O�f<N`U�C�.�
W�P��@9`5��[O_1MתL�7C�XC��`�R�m����P�h��=Y&<����A�N�ʘq���>| K��cܸ���R����t!To�����:Z��?���(eB��2O�f�Tg)`�Vt��bYEZ�����V���*)9�wew�*`���%��צ6���X] �ۄb�y>�l�8:��S�ʡΜA��ݯ~
w��e�Z��FT�v��!y�:x+y��[Ά�q# �?���2����=q����N���'$�ًr��cs���{�H��D�/����%a<O���%���H5=B��]�>�a2_���/�|���
����/�J��Pa0��{��u�!��*��I��rY����݋�l�	�3 -��]�x�U��ژ��2ﲨ�fwߠW�_Z�����e@��4�� ���ASfx���V�Q�l�L��� t��MHWo@�� d�P�
R��%u��bz�C%DC�s2�E��c��^y]=�iO�t��@�J��Fcp��po6��� o�uT�xEUGrE�t}5�ᑊ�w�
�<z�Is��ک��S�K�Z���L���%���NRլ�d�El���kҢ� ��s@t����g�Xs7���{�o�y����������r�c�$$��4m�yF�K7���s�Җ~t�����9$��س�i ����U�V����ku%�{?&��m�`�/�e	�π�����!�h����G`7=��g��`"A�c7��>�>"Q32y]m�.t�=���ш�<"�F�T	=$��3�R��zeN`m"���y 惾z�/AN,_Y���O��i$��g|�%�k_�xp5 su����e�{#&����Bjc}���ؙD�	n`6�Ej�u��S/)�S����?}E&w��3���Un��������/�_m��D2�v3��������n����hnJ��H5n��M�9��0K���}i�!qP���r�w�[;�K1�ا�2�	�
%K��9��N��)5�e���>7�R�ԄxYv�H�\����	�l{���z� zݩ ʯ��yJ�e	�9��9i;�_��N	�@g�QV�K+�^�o\�P@^:K�2�z��)s� ��Ò��3"Ƭ���M�" '���"݇G���}��{X�l�;��'.P���f'nӊ?J��zN�`3��pq7{��4�ѽ����Qg�N�P��j���I<�q�7�H�y5����������x�xf.�4����T#̚P&���;a2�p���vW��g5ㅐu?4�U����-�ߦ}\�D�>�#]�#�����ȃ�7A��\MR�|�n4����~�{X�qz�J��!Ot����3$Wѿ��]�Nkۻ���O?%W<x��@$�-���ğ�F{~V�Sy��/�R
|�7��'%�{�4@�8��1���
U�����b{$���&rl8�����e��r�P]�DX���Y-��Z2:]
�u��ixc����U�"�e���� rnPًQ/�6�x�d�xk���5)�*>���A�p�1u�#@O�%���6�OIRo��9�t0,�]�R�.ڿ3��uI�6�ݛ�C<萶����]`}ς�׋O���	Kp�|�pj�g�r|��ʱ꯾��a�8|���S�E��o�zR�-��ҋ�:=�!5t�.����(PH k�)�߱�t�:\���㷃���)�
D��x<I^ϛ	�ߝ��|�����Z��fq��[��Q�&Z���/l��Ԟ=�>��}�y��=߆�'�e���%_��DT�����P��?�D��m�ӻ/��������!��^���A�� ʛ;��B����?t��v	����j\J.i�T^��Y�D�
Vȅ�=@V�&��C�'蛖W��ra��[�{����&,��=�����e�F#��r}"#�.���z��\���{,'���Ꟛ�َ#�j�[#�GS��L�p⸻�=�J0��C�}2�����l�)	�~Rڔ'����1;��f�ׁe$M�!*���+�m���V���2,w���^ۿ c���x�,{y�egN"�` E4`�qy:$���"�:xj�Q$6_�&�M�q+q�/D8�O���c�޷5\yt2]��^�d\�T06��+%�fs�� ��瀲js2�KR���|�I�>���j�v�����Ɉ�EeF0%�3�B[�(��1�"&Y���Gݱ�,��g�����q��?���Gӳ��Ĭo�&��}>a��}D���gI��
':�26|^=��_�=~�`�Ch:��*��x �DL����܈�$��w�Ω����"���E�$��]�n��!+[=G�	����	'��xQ@H�-Yl���Y`�0�\�6�Zl8�k�$t��oV�Y(^��!ꫮ�Ԏ�eVu��̃�u-�UPR�Ўq/��[�r��ɽ�vm�-(rt�*ݦc��a��t�!�+WEr*��U�IM�)�]�X1���#W G�W����4����[X�����U/ Rܤni��?�!zM)m +�_+P&=k�G��g/�βd䗒'���O��>�=\��^b�h�b���e+\uF���a��Ú��� h�Q�
gm��'�ƍ��W�&����	��O4�e����="<{S�'��e��{������r|x\�	� U��v��>�WӞ�0����cc�?�I�-5�#������ic勄yw�w��aI"�l��e`,a�!Q{������i��y���Mxt�p�~+���{_�Epf��萄�u�O�fۈ�fw�9��,�֡B�P�0���bݜ ���\��e�I-�M�ǪA"�^8:�!�%�����t!2H�?���w2BFz�7<��H'+ۛ�)Ӛ��:���?�j���y�V��sG�K��:���\��V���8�OLe ���C Ԗڝm�<9|��G���?Ĩ��,��Sa��x�i�Y�-�k�<h��5?��#��<12s҈:hQ]l�m�A�M��ų���^Y@jQ.a��W*r#�bH����qT's+}ל�n��.��'��#����U>��?�dG�]��)����j➃ħl�=��;��+!�0�����Ƈ���	9@���~�h>W_�,7���/NL`}~�Sx���в�-W�G U(K�^;!��ꃃr���>K�g��OC����T��EÓ���I}�G��(��!��f��Q4@���!8S�/���*�����47�<B��ܻ���s0�^-'�rA`�m��Sh0�G�Jzۈ���	=&����2�}�!d��永�-��S�w���6���rc��9��y�(��h�8�
�҆�&h������ʱ�n*`g�ٖCbM����~B�:�?�ⓧ��Y������q����T������rF�����p�@�w���q��9�&��JZ��$q�y��@��x���ӷOH3��-`
��@�9�8��8K��r�<�F�F�`q�7ͦ���bqӅxI��!�\�C)WF�du�&B˰�ە����
���Nȹj���c&H���9p�o���2�:`�h��#O��`���(Ҟ�x&#��Y�?*��b�O�PZn�n�W �px�����z��_�*12u� �X'�?�V��3�V��W>���O�"<��="M���v��r��H!��5:��!*��GMtya�z�(_���簂c����Q�R�t��#�����k}�B���������7�|�;��veG�W ��i��~u������&>����<��2��`���f�$�:e�s�#�'�;��$�=�~�l#Ⳟ�DH<B�@Q�M�9�܁��ń���O�Up�=��Gz+�$9�v��W^I ���m�?�,O���q�����5f,�r�S@�g�7(�N`�>/��]k�f�!����{���L��͝a��U��>d�B,�7�l �
�Q�T�Q�z6�� ��%/$���h��<�İ��=��-�%�@�r�;T�'��\w3~��F����b�v�"�+Y�F0�]O����G�Q9���4���n�5J�<��<TeW��M�n�`~��+�@�"��!��#��⺗�hD�:�m�������R�&�V�R��˩޲y�&��pT��*�ʘݍ�#_�iZ�з�VJq8'B��ssM�#-lvB�n��0��~
!���;Z�Kְkob��4m�>���yq��+y��ɎT�s�9�y���j��.��L�)P���~�2o$/U|DPPƬ���R�6�m-�q]��^��Cby�An��"�P�(Ht&zd�5�wB�v�α~B�R��rg�D�����ـ+~��x�Q*���Q��9UJ9��/�E�ФVj��WOo�[O)����+�E�����ޒ�{��}�N@���|m��|+�Nl�*�q�KX�Z�a�/�<$��?�Ek�l���E��R\8�_���c��}H"|U�~��1���h"+1<s�P,�2�c�Q���<�B�|f`���~��N=��Q�������!A)Eʳ�~�~���Agr�s�;��8Q����q��]`*��d��#�k>�6���0�Ѥ�_©ٯ�9�J�-Lz��oQ�q��/�a0HP�i����!���>���s��S�&�3��~k���3����%�X1��{ߘ��t�N�b{v�-ZO����n���~��=X0�G�Ք�i:��F��\V9�Y�c]��#��O����ђC���#�Ì]UK.�Uܫ*�w�����7gѕ�*�5L,m3��b�Ӳl���vh���P>�Xz��գ�8�\f'�@�nt8��?�-�Ŗ۷GU(�p�:��[���Z6�Eiޖ⾘�o���8X�g��5-��1���>��"i���Jy��������N�RAēƖ�w�k3��L�� q��M>�_lvS�TU]1�櫎��DM	���P�aT���T�N�^'�>�{�}%��¹��b���H%p�mu�_��V
忠�XI��iC�F�Om�hf��J���^�x�y�������'���55���_iH�%..�d��Wd��!���_/�/��G.�[Ku��#��.�t�A9#���/�Hg�Xx�����w!֧�Ex�P.���Tet:+B�[0G�r(��/%N1�z���Z����B��w����,-g��̜�������2��
\��"�{�`�3�2�&�X��ap���*�j�p0����|h���D>��ј4�qw�~&���~_���;���.�_��������/�bh�l[=��o,h�%@|���w�ԧ�� D5�J���s��%WT�5�2�6��������/�Io�^xRmX'_�c��6��~���+���MXR	ܤ��\OI��D��_}kcc`��`�����X7G�-����J.��^g<���rsoNs�T��Y��A�5kGk�ȍ���I_���b��ѱ��T�Z�˓��wڣ��xJ�(޸SB�<Gg�=m��q)Z8.?##��K& |J���Fֵ����DRL� h�̚��t`������#]ޠ%��_�$�ߒ��g@R�X�tpT����������$�'�Ha@�ʣ�xT�~���WY�t.�#�2+"wa�Zpkmkܤ�������Z>l��ŭ��ZYld��P�U�;�6�L�ߘawiK�s;[;�#�����1�t�OG"*�8=?z�@���*�$����Ar"9*f��o�����꼼Nh���xMAs 0o��w(OUU�j�kp�N�`{�k����c4�D#���@�j���������.��So���b-�t�a{Hx�r�Q�$����O��h�b�w�%��	��Z�����{�����û�8���2T��pi%^vN���d�m7ꥨ �����ҏa��	���}%&��ە�� Ͱ����nKIgoV �u)��f3�%P~ҫr��>ڊ��������Q�l1O�f��b�q*���%�P��Nu��&�����JB�0����	,��>뽍�E���%�'�T:�w?RV���Վgv�Y$�d���ǭ���uM
���?7��T�4P���sh�t�ǡ�gsT������Ǟ��
�^n2�3F$!S�7ߌ;n��G���ӌ3W�[����-�K/�wE�42&�<gQީ�+R~w����dk��{2�p�<;�x�t�?'�@v�:�K�\��ɅAC�Jb�a�OۂW��_�J�]�NG�9��l'M�)��TH�6����xe�`�W����D�a(n��w��ӌj_�p)ә�/�����c�ET��^�۽��x1�֕��!,Mz�@�6��X���
���Yݜ��T�������{�e���-"��];O��/FrD+�,Y`$߁���R>o��X�h����;e�X�` �l�!�l�7I;IZTHqm����Im~�z���C��"-h�f�wX�}�S���M�?�_���ɗ_��	�|f��;�f�Q���H��Hb�/lݱ�Mn��V�8����MpI̍�y��� �&)�mV�UG�3o�M�3m����C�"����!���}mWx.~ze�sC���<�D�X�E�$;��|��9��q��9�����L������-�JS���f�E������!q��o�࣊��֦�P���1���U�\�? R�P���8��K���\��)R�rRx��Fj9�@LV�*��{���X*��W��^M.S=�@��q�F�Ua����Y�^1�}����k���2�o�B${��GLn"
���kk@"�vK��ԏ�GLp"���'�V%����v��WW� �J�@Z�֩&֌%$X� �TQ<$�~>ΡK���M��R[���u��1B&+*z�Urv�SZ/2�A<�5ki��Rx�Pb��P�{��Me+s΅[���B����̟������I6|͐��L]��<�-L���-�ӽ�g�E��Ҹ�ؽB�<�lq��Q��x��POE�C�Nc~�b·f|��l^���W��5�(MA�M[D����@Y�r�����8ҝ^	r7U�7���bPl���3��
�`݃�����E\�T h�'�_8�-Y��2^�{����|bޓbt7�̬%��m�fi����5٢ݗ混#��1v˴d�S��J@�3*pDM{�|�$$x���ǀ�<�v��Y�࿠�5@�,{��r�ל�t� �� ��g�vm���>^m"[��k���T���3���+	�{̄&eR��U��k���j\�{�b_5p�	K�wbOn@��u���mv��T����6�����:"D��!:3��k�W�qP��Q��vǊ�v	�f�����E��Q?�:<���W��Ր���E�Њ��\]K�Ɩ�P�U�.?W�)�]4{1$�|��u�0.�����(�}����R�'@���uX���y�>,g%�rc��(�c�I0'~�n���$2�)�V"U:<�޼��Q�L���*N�9<��ԑ;ӀU��a�<�ww�Zl�|�-��e8��Tk�a�kv����&0��	ǫ�:pa)�ٲ��$����ؘ��+X�'���E��%��ߚv8�,��@b V7�'�{��vL��B�����U��i�N�"̵�4*�c��4H�*�?b��d�<sa� u=^���xj��rj�
�$���U5�b�4��L����y�-�7*E�[���� �O���M�������L=�0���TC	�D<o-�[vւ�����C�]�,�P[pP���ϐN�1�C�u�3�� =����{l�%��=�C�*
��Ű_��,��,�d`0�������g�#���-��:�R�t�&x���ۋ=��A��v�{�dP�]�>�T��<ø��S� jq�p'����T����u�	ő;�8B�aTa'A���R�����0�/Ȋ��Se>��{B|��ϵ�&`A�L�������l���#ʺ�N�k7�6m����z�f8�,��AL0�a ɋ�q��cU���z�j_�(oຣMF]���	��>�@�(�ò�#:4�P4s#|�:�bx�ft(u}�\��{�w���US����.���R%~�uk:d�㚲���������N]JE��D����`���$��	��[i,�,�QV/x
��O{�(��D�/�Qv�IG��i����?)��h��R�O,,��?��>��"�x0t{���޶H�"��B��<r�;����J���{�m�ލ#ee[cp�CWɶ|W^��C�����.�E�`"t#A��]�8��K���F���xh��(��	�f��O>�lih��RfS�~�z�W<��rO���/��=������X2IQ��,�wj����1����I�sf1u/�����
��X,��$
�T���;��u���� 4c����:ZK��W��C��`<Լ��&~�ƤI�oh�^��'#�?��ټz�QB�H�R�@1���0�/{Z7��ؤl���ὅ�A(2�ƸXmh�,�E"cS�i���9OTy�6@��g|�"�yMp����j֩�+��@���>�����n2��nĿ�E��e���-sB�o�F�sI(hi> Rs�����T�(��gq��>)x(�s�������6���S#��8d���xN9�n1{�t�d����w��]vemSY�:�T��hd ���m�x�qq/J��P���7
q��z�ߒ�2�&�{�,�b?{z��� �ސ�ںGn&��-�b�O4c��H�e����i��<1	�x�x�0�ub�\=K����7�2~$8����dN�+X��]Z��v�8Л[��$���<YP�;�C.��o��{f=
��X,��[;����S4ہ(���Z~�˼3ф�D4Q�Gk�^y���;/aյ�zJ\J���v�+�t*|���e���g�i������3t"�go/�jp��1�}��/~��&͞��J�,H$V��@$�� ����iWg��*�5��h�s�
]�j[���|����# T���+~�O���J���8 �pm��:�H��\U*ǙQDp���f�<Dk��F�0N��p��-���3� �|Q�	�T�C�ޭ�K�@`D��r����Ч���/�eWW( t�{���-���S䴨�_?q������lV��v��K��M���La�^��L%�Q�L����C�&)ݞ2����ȳg�\�DC��2��Le5�'ڄ��8c��1��N��P��䱬v�#����(�Y���g����� �_�hO��5R�F��
��ζ.���=�̀U~'|�s#ԩ��YZR:�~�h��;�-��RJ�������=h�����_��X�����?w��n}���{��$�@����̀#�zӰ�=��P�Z�&��ʄ
;X������6�^!�v,֎��4�/�7lF��͆�C�?���H�ͼ1����JU���O���X}�Vm��V�\�&V-`F��6��&���N�3j����4�ӽAJ��'� eC�	\�&��sXS���Qc5��2�X��D�J�����ΐ0�JK�f�^�c݀<a99P�O{qX���j�Ԋ-B�DF�4[H�Ul�t���+���_DE�~���B�UN�����4�9a���l������l^��ڔ�r�-ß>�|���vHq�kU0d5�䱥�0�������?���;�k��G�������g��^A"�GI�yЩ�O �~��G��hUTb�:DMӱNkM9 �f��&:1I'P��hX5h��7��;�x�fgFȑr�J��m���N,û��s7�I�
�M��s3���.t
ٳ"�dy0+�z~_�r�5D8y��j��	6�twAi�l$wo�mG\&�h�V<�׳��w`�5��<�~D�w1��W2�zo�|�
��v���٢��	��`��.�\��|i�P��;�:�`ɽ���6B�	b���<����e6����L5�'ȩ��ކ��aH�ٍ#�($5v/�ҵpY~3*����]�U���0��{�t��Ō`f�X!��G�Oå��^�a�@��*蔜~}��i��w�J�F9lW�6�O
� ǿ-�okse�e/���� /�-:��vI���
qQmB�H�TߖI��o�$Y��V��ڣ@��ѿp0��nz#���?�2h\�C�x�wfqئs�@3P�x���C��mg��¾O]a�:��_�~~� X��q=�'�b�±~@xg6����/�͒��`�<��2磕_+XzpyQ�WTGz��?�y��+v�	kDLe�]�豝��f�aL�8��/סO�G8g���g��9{�}[PVX�9y�Zr+�����nKK'k����j�	�4�2\��$F�a0�J@��2�d�:�|���5H�vt�jsO,kqyI��͈4�3o���>Ƽ����K�����ʛ8��N�
R�� ��g>JD��[�����-u��$\�9G7|�_%&p�k�64��";� i�;�v�F���BIy�3[�un��'�@$����Z��\��r�~���a�^�CeP�ALL��@Շ}L�׹rSKC�݃t�
��hj%��Z�5��%?�f��Vs������ 2���0������m9x;u��]��P�,��U����ѤW��3��-�+�v�xG��p]eI"����ׄR论=-�.5JKt��ɾW�Q�96^�t/.��N��"+Cz�>�Հ�&��$r莓�v_Q1>���f)�(�unq�@kl�x�mZ�^`8��f�~�;���^I���p*ݱ���^
�H0lyΑI�6��8
p���vp3�;���֕<[�$�}62� /�>��ή�>��z���=�dy���
���grR���KY�A��j﨎d�f���#h�R�������3m�>I������Mh�r��~J���O=�1��i��*����3������#���Q�5v�2�O<Q�� IѼz3 ��[�؉X?��PJ^aE��<{�������I?����x�'.�G���3175l�L�ll�_徿꣸�+ᛡ�<�b	���Q��wHNX6Ɏ��~�_ ���E'T�.�����P�vL�ja��u���*]�q�vA^����>M����b?��U�W��-&j\�kTg����Z��(��W �rR�UǺt�w����G
�v�7��|Ⱥ3(!��	�|�&�+Z&���
ìW�Y��|W����fB���!.�p�/Y���5ik�2k< �l����]������U��h�+�Ǘ��H�������OH�h�M�������'�U�eő���3�V�m�Ҙ�y���9A�=]̈_�}�!��0��l��/ӵ9�cU#I��x
�G����L9��k��x���V�f�C��} $���<(�̢'6g뱺�Q��9�tϘa�l��2(X|��Q�=��Q��P�=�|�xҿ'������(���Hی�l��īs�o*�ҕAUOչ��=ۥ�0:�(0|\с�	�R��3}nҰ��U[ ��0) zL��!f�|~���Zq�k��J��� �Z�݁��ak�a}�5XxC��<X뻗����O��|����Ed���L�|��ّ�[�ϐJ�M��nO�gEFi��{ ;t4�eJ��Z���|����ݟ�M��K)'v�#����ܸP�y������Q��m���FG�ߵP{C
���"?x{qKIN�mpV�b5��t'&�6e���K^M�B�v­)��@t#���8@�o:�c� �E�I�p��(��:��}���!֌��6��N���8D�P;�;
�c��i�J��d5L�Y�����8��'�GE�n�s���k�$�b�A�281��|��3"Ȳ+'6��{�l���,�f�D	���O&�M$4G8�ʫ��ziꡁ����ͦ3����B/S�1��KxR�29����Q%����ȑs�����]�Г�|�uM��V gSl�����,��7W��P����Θ�c9L�PUl�8���F&�G�n?=4!zI�F�K�Hgy+)2�f���Y;hA^>�"]\>�hO���m��I5����N�m����2���
6E�K��ݬ��]�f�"*�,�C'�C
�5)T�����a��k�d&�,�����U]�	���!���Q��v����._����X�N�]1���l��0(z�JA���\��W��_o�,׻f�R�����z#m�=�F�bX_����@k�ԃ��-��C��%[��W��}�"x ��A<���F��z�QX��hp3�O�ZM@y��*�����z���<��Afb�r\��%��?&����z�HnU�q�&�+hW�/5b�9����Eص߬���6rj.Vc���/���r��<~�}kT=���:g�ĉ�2gos�"X-U�U��&��t�O�yW�f�	5�C�&� eDK�O��	LK�*"Ve�Tᱨ#ί}��k>�������T윆c�Bgf�1MxD��
�O��o0s��"���Kt�]TA-P��Z��2��?�����"A�np��TFAn�I<h�:)�}��I6ߊ�� �Yx
�lJa:bU�	�$b�ek%��C/�kT�P�e��L�g��=��i(>���SQ:[ ��a�-�n�{L�����jۊ�g�C�=SR��T��CI�_�����0uo��2�0�l~����xpM[�ջ��gK�ɷ;|V�[���x�v���� �پ�=�ܴG�I-1�`\����vLr�#COs��095�gr�x��t�æ���x�A���&�٠b[�xvIn��0߮<��q�m>Ãu�8��?=�m��DT�H�K��$��	���m�V�|��	�'.I���'ɵx��z�C�:|wc�.}������w�q�����}�W���Rv^�Ϸ��4����a���������6�P�e���y&:i判�a�Hh#�r���;܍�\�Bƛc��n������7�`����r`�	������6U�9w����И����D�f{��}OBw�ۨ���ELy�}�?��v�I��@by(��.HL����� �Nt�V�}"��n"���� ��v�+�NG�C��?afxx�6�����ڥ%211gR�@-r�ŋ�.i|O���o��\R�Ƀ��4�J��%����R��½]V���N��Ӄ:�����䆍^��0n�Wt�> W�����Z���S���+�?�E$0%�3E�Ȯ[��-�T"��E�Bb9�vP��Y�=�y�����	T>V�(FAb��*�B�J�ٖ��=��Uk����*�gޠ&L\��_2�d�����{9����(wN�������}^I�n{:�R
�B6�H�z�s��4� \�S9�x6L��m�k����?답=Bo�K(�b7X�_2���@��H� �8I]�ckaAE��[��C~$�^P��؏U������:�g����G�)/9�;�W0#!�.~�㖧;s�f���������#.Y��K)qIo�w�B�s!a�+@-�߆Y�w����*by���z��CUKad�fa�d��IP�*����!^���~x�P j�\��J���^��~D��Q�P�=�`aA�(��WqG@��Z剙[��c���v'����tL�P�.��� ������Q�T
B7, ��Бgyh��СfIv���������Z�ܓh�_|�s�מ�)I귵�K�������!�\�~�z~GX��XR܏-����c��T�+,�x�����q���)6R�%qL,��A��a�U��6�mq	v3��q��`(dB�bq�@$L�t���Ӵ���}��H��'�������eCN���0��E2��z/i�շ��
�:�q�������k|͗�Z03���k�R\�GA9M�x����@Ec �1h�Rh�5feE��JpO��#��7F��[���ӓ�[�
1�|��V++ߠ�`S������E��á��x��@eTzf65���BT�*������!���E���[d'���y(0�w���8M�7�1��T�>���@[k�@X���v���n��/$�C�D,i���T~j��i%p<'�mj��~���_@�s�G;7�cq6� > T>���w5`,�*u�#t�>�5[3�7�E=��z�UTLofw-0�.�ϱV^�`��A�L2���N� ��o�ü�A�=���"c�;�X-����;S��5�A�1h��@�(_7�";6�u470�L�4����\J�u r �i3�Ǎ��jxT�I���m�Wf .��6z���tC�8b'�����Pm~� ��bˊ�`�#,_@��o���%�n��naD>MT������g{(����1��R�e�y�VT��Cv'���㮷@�H~�s�����Z�6�.Ģ��*s�"?BZ5�|.�a�P���6������T�s�y�m�J���u���:�rO}40S�J��FJ�iX`���u6^��~GS���������_4�7R&�ѭ��S�Srs[Ez�I�n%7%%���N��@�,���W�-
;�Nԅ+�Փ��Sx����?�P�
��
U�]�ltM�DfB?kд�8?����\gx@�Įq����iN� #��,��Rѷzu�x!2&r�*<��o�ײ��e��Z�a��bS`��c?���N@����{��p*�d�����'\pX��hl��7?�dtW�j��rb�� |�9�{�N�9���Y�@�˰��-`t{����I_VZT�@2K�LϤxI�wȴOG�&�u���Ϥ���ϗ�@K��n��&��z;����`����%悩�� ǌ�����Cu~C���^��R.�-?h��K
~,�����+upx@�i������0�.���B'��Ӝ^�2��j*_e^�x�D�+"���h�oޱ"���7�����Ԋ��,�)[,K4�T �c��� �} �G�W6ۢ��<�L��X���T���eԂ��+�5��Jw&-֠���ͻ��@�硷̐s�:P�@-�Tʵ����U��oͣ+*��!����I� ��7}�T�g��^�ؽDX�E2E�6	/�ؐE{�fH��[7������H�������¦x�xC4���`��W�ҍw�+�<��i�<�Y�")?����k��)��b�O;�8����Y�����Y���E ���䄋�c�^��d��i8��=Ŕxň�����i$fN����b�� ʭ�ˡl0�|L������C� ��t�����ބ-�:�UeA�I�ZM@2?l�Z�ju�����e����+˶^��ҽ�����/�"l[��'�p��O�7yo�-�ٌ+��骋Kgs�ʄ�3�Xl
5_�eB.�������^tu��$�]R�S�Kxh��#KW��6����i�<M>�ⷢ��i���'������Ø�#����_�!Q�o��SLG�^҂�~�,���StC�;З�7-�3�*�@S�ͽ>��l�MO�R|}r@�݋c���G��KE�U��,�����+�
�����z��"wf�nI�H�o�i+`��Nr��ݍ����R��Q��y�Y��Q,�I��r��$�L��T��8���ߏ����WU�[s����5����:��]#`�k���KL�W
w
�-$��ك�����U1�^�6�K����t䛩�]uV6
���f�8'G�LO5��U�Y�bN�Տ2/��Jt4w�pv�l�!X�niK'v�N5ѽ*��r����Wh0S�%8J�$��>"�$X��Ȼ���:hAG�0�W��?EJ�i�~�m8|�)� LK���V�_\���zl4ϐ��,	�ղ��b���L�	_ə}��^�e�?����=P�j��r�*�34pw}�t�%�Px�a�G�s��O滇���o/��W�TŅ�*:Y����4��90zdC��fȄ$p(]�1f�S�4R��[@_������^ ����C5�u��Ц�������o��
c�W?x_��E��H���n��59-q���Q �Iw�a�-�����p|�OP�?R��۔���~����Y1òx*1A�q�>��֦hZט˽s�7}n�l��(/M�D�t=[c[��6W�hk�/�ΗO�I2����9�\�*5��y��j�C^3�:O�� U!格���@0� ���������s^��n_�I�<��Ǯq�� 8�]f�{�����Z��V��8n�q�r���_k���ݤ��P�+Y�$����q��E)���)U�r�2���m��y��&͝T9������R���+sl BHd �A�3���;Y<�B)+�7��Pȭ��@2LQ���8~Y8�.]�����;�K�v�9�����Ԣv��3-��@<�c�:���E��&a:*|��q��p0Qu�h�G��f����Y�d��UH咻��@w��qi�� yq�6�"�k�T������9%:��� J�[a^T�2Zo4�O��x��Ճ=،.�[�oT-�����p�4�<3Aߏ	��^u�1�B�ɉ����:ضdG��x'3b��'"�ZV���$��8���,� �`jܭ�@��Qf�����녾�AS`��k$#��$�f���̫1J~�ot�S���?)t��T+��o�v����$ ��Ó��杴��ٞ�J���I�?�����[�b��i򟳳�t�K��h�_d&}��YlRN`�����:/��wk'��Q��q���A;u�Q��MML�7]b6$}��/|�Ŧ�=��}QO�^�$Ǟ>e�gxN:w�ћ_s\�@��}��@ېy��`���=5�n��ڝ��W�]��H%��GE|��Y�\Oe��,���½{�(��N�A�0bη'�$���?��dH�e�h�gH��Kzi<؝Y9v�T��O�!�@�{�� n�Dz�&=���N��n��Cq��^���RJza�4ߜj��,)O�v=�+�_��Mv0�tT�w%Zd+�SG@�f#5xR����kY�så.��/��Q��T�z]ޣ����=R�NA�R���(N����.����"���}N�VL�O���/zẏ��D�-�Tb��
��"��S�v+�#|+&(�oEP�DOw�����4o�~���ūM������%�!G�0�A��_c�b�
�ϥ�[���@o�h�ht]mD�:HN����]�=n3�+T�K���AS���|���0�≯�-g��?���yD��9�pzlW����n"�`.����5�a����_q3�J���f0�n7�LO��Lׄ>�(]��~��� �p�G-=2!˱*c�H�I�c�SU����*�f0�p2-V-Ac%��O�J����� ��ũ���0�!<�p�e���Ѥ�9�7�ePv�:^RL��lW�[ͯ-qC���/|]sVWt�_N�M�9NV�2@ϡ{M��<�E�K���r��=QM1'��ʨ:����ȹL0�k�C�en>�#��]���K2��%���QYڄxtҮ�� ����٥���9?��tk���Q�|޼��@��J��E��K��nc�	ʥ
��;.eU����X�$���~�����N����$]L��c�l�Ϟ�P��,�1|�t~_
5K|Cn�6e���X�?er����5J���0�-h:#7$bq�G�lV�vA<dU�|]��H��� w�X<��sµ���;SJ�s�ܲ�Ǧ�aP���Ԙ�q�h}G���f�,����#�������Z�V@W9T�����ĩ�qrj64;Z�w�m�.����vG�^��2v��$u%����NN�8����@$UES�}�|��7�>fL��أ�u�Ԏ�0'D�=Lb��������|���B�<e���
�~ڊZ�f��'��3�[ǃ�x�(�a���U�I}�$H@�,��; 8�~�4<D��'I4}�D6h��K����]ۯ���X;١��`\{��QBp����-�ULO��p�A�����ܭ?��;cQ,IA�"F�ڴ�wWC��1����/@�E��R���#m"c�";�n�AڤD�\T:a�<�J�����>�a��a)g��o��sQ�[xv��M�r���B�|��cm�N;�(��@=J�a�2�;��P a�O�/��tw���o~w��K�њ���/�]�hB�H��U��._��~�Ҧ�>�kgo����#p��%RAŤ�j|����B�||�ƴ=��<�HRc���)������7'�$�����yN%����z�Ӆ���qK v����B��̙VwY0�4#�(�\��X�f�`�����YoC�iiэ�%6�ڨo&�5�W
��n���LP6���O���UW�#�4-���G��]Ly8�S�'�!�R=�ܻ*r��Q����Ֆ��0\��P�Ǉ.�y���̱�~�=%?܆�Z�[r����@�[^oy�3rw��ٙ驁�3������QL��1�+�#u�w>�k:��E��}����*-��oK/�H,�"`ܯ��.;_�>��R�+3e���Z�)�|�5�FD6�J�#��UQ`�3�9�ɸ�������_adt�����s���*�����eU�݂���O�AFS��ӌx鼌�x?lԾ�eu{�K��P��ա{�Q��h�8�G��;�W;�	���·f�5�f	^a���W1i��=%k�
p��߆a�?bZ���Bm���o��lw5t���u�-���#����^:~�O�dzs_��
����4$T(��g|t�b�zi��r�٦���}�1�3��	����4�R��X�x%��ҽV�)�ΧF�s�5fL`�c4߁�ٸ��(Fe�������s+�>Ii���M������4�a���ӓ�d�颙�u�P��6�>��m�X���ps���D�k������|��ܚ������^��,�^ix�#
H�}�þ����+��1�1�@�� �t5\�Զz;f��C�hc�z�џ�H�2��ĹM��8}��T� \��M�*�
�u�����Ҏ[>D�b��!�V�weM{58Q4�U�����]��r6V�J�(�QuQ.y�4�Lv�}S����+{h� �<�-G*J
�>�o�;~�~��0 �OSx���4�"��G�.�I�r��Ҷ��ح*���v{o���]�1`+��wz�2���{��pE3�rq��e�����v%�*><:i%�F�Y.�s��������}�\�F�ky>S��E1P^[�*�q���ʗcXl�����[F�I�>U3��<t�=��Y�ш�=m�
ƅ�A+����6yӤ<^���<��M�ѐޗ>Hi��w�+�R{�2��諄~wu���t@q:�X-y�>+5PD���f Z�D���.�ew�o��<Z�i��&^{D'�G�œ�3�-)��2s#v����C�F+.R��oa%{2�pE���<��J��Ŧ����ұ!��7�Z_�&78˿�G2�$�n�~�Tq�sS�?�A�*�Y��ɔ��[�6]tE�$%V�-���a�.Z�M;rE�.��Uqڕ(��9���$V�z�h��'���]e�g�vT�jP/��AP��$�53�����qQ�|�-/�]�?Y�0�l����ޢ�ciX�>ƄP(�q#i�U����#�� )���Ce���X�e�2,�/��;=df	���,N�J���Е��KO⏸[Ã�EGߙ�3��;��hk4,6q/��\bL{��G��K��J��2��ݕ.^'���1�I%V��6o~���p�=��n^��뼟Z&79
���?�wm���ǯ�>غ��k�;*���ѐ*�E,A��A;A�y
G|K�
��Y*M�hϗ��B�9�왍���n�W�M��Jw�
�h�ZN�	�[բ�N�;�ͬre��>l;)�E(>90B�K^�b�_�J�覼�O��z9��{������%��}�F��D����&zW�N��.ƹ*m-X��lz�����,iuj��b��?��k; c� 3C%Ϙb���ĭ@�K�p׿&��II/q"F�C�{I47º(|����(�)�fD-]O�K���jY�Y����x�*0)�ɜ�[k\��?,(<�mwo`%�"��̈́��{��|ˎ:��:n^�W���BH��Iu�����1�ua���<<t5�VذǪ�H]����VȺ��M���Y_�bJ������B�2B%u*v�e���v[�~���;���l���8���i�����dS�?G)T�iH��
�ʱj��^�b	+]�3x|2z�)� �]�!r�޵�2��&d�tW�c��@�<���L��Kq۵��b�|�h>޲�r�&�BF��c��F�(�O�+��|�]EK�콐�l�WOS�D�M��H�Y#* /����,�[����(����Y��$K�{�"�m:ٟ����:L�vy�PC�lP��Vk�E��l�����C�@�&0A���JO�G�ye��e���X�G.c��@Z(z`�3v����t2���!����I�tѲ(��#~� z�c'=����\��\~6���������v:������ޕ����F*E�������&pّ���� ��QE���}�A����@p<�����-ٟmj�9��7N9p7��=�~��iQm���H�Ck�K��'8�X����� n*�6@�e
��uKͪ}b��	䌋泓���A{�0�5��\j�j�D�:Q����%m����-��1�Q���_�f���ӈ��@�e3�@uN;�5�b`cd�;�Ӓ�V�B�y76W)���0�J��Ғ��f)Z7;�|J���j/���gTۋ�.Bѿ,��/�6������}Li��$��ѥ�cO>�:oU(4:~Q���x�o��	��l
��C%&�\����:��ގjM]����ElIho������nE����ٛ�J���q/)�fʢ�GM2�K	f�����H�p����c�Ne�~�KLC�]w�pyr,&��:j��	�ԡ�q��S�۵��J�>�FΤ�����P�U�Ԟ�D���n���^�ĝeh��h����:�EQ�z����r^�L�ً�D��RJ�-��,n�@�3`�V�6�\F���.����8P�F�,=:XV��`9a�1�ꗑ����;*W�F�_�������a��ݴ�BHrt�!X�'�&­�7|tN|xĜŷ�X�=%���Lp)�+Ɛ����ԩ K
}Q�t�~iPZ��Τ7NLLj:�R�ӂZ$�"�Q��FoEJ�b�(��,�k����_j�E�<���كb 7��CR��5<����drD��[�(}TC��1��b�(�kW�ʜH-�:EF�m<�'�9�MIĜ4}<<��׆�}�$_w7"�8�7ۀ��$J��_��E�w�..季"�|�`N@X��.�:껌���B֫����E��!�CY���9D��j�Z��g٧P$�Ct�E��M�lm��
=����9m=e^����;TS"��O���j< ����k�lv��g���w�)���	�Y'e��k6��)G�3e��q�|�K�+0(�Y��D�I��Id>�[��F5�A��-m�Ş*��7w�F�hdg��o�� G��2H>��lL}��������R�U�����һC�n����[�+���	|�+�F�Z�Ǣ��
s�dr-�����X��35?�>0���u�C������l��da�̸���#C)�	m���u��t ��Ү(���������
�}��U9)�����W�*����ۇ5AEg��J��/ �����ջ��˕A1Ɩ_�7�qk�j������5(y��4t˵'�Un�r3�t����z����J�)Io#��] �H�c�'�yòy%tw���Y`�(���9�$�jE��y�za�Zib�8H���1's�ǧ�o�%7��t������s�O�A�*^j�A�S'�/b�v�7(_����7I�~�F�X��-�R��d?�D����5yn� ��o��ݴL�2c�a,�$챌�O���R�3�7�f���9�[��|��C?|�%ߪm���t-b_�@]Qk��c�p����	�:�7/?�h6��&15���y0'qXϦ�koz�"�L��Y�ɫ&���@'���S�֌�9z�S�D,RÌ����6��bm5�V}��"`�A��h)�)��r��z9�cha�%=�^�	/�g���k��~ُ����#:����l��n�NΫ���$%�#��O�Z,�$k��4�XZ��#@3UdW N"@_�Uz�����ٝ��n:Ϩ3P?���6a�W9�	��2��ƞMn�r�a�v��ɒ��̽�3Ӯu5��X��V۰�A&b�|Yv�C�
�%�&y�3����
��[����p����ڀn�.��\���D`1��Ys�`@��X���ߦ5>ɋ8��ˇ���N�̞�ݭ�\g��8�X"�;��d�w�:%��VYZM��
�!0r�Y�� T&�Sm;�W[�26�"ĹSq��}l>���f�\�Q<f̴M�Y��'��Y�p$�*-%��D���*�ڬ�/r�8�Y���ȗ��J�����P��*N�Ta؅&���r���O�s���VyH�=	<m<�U�"�[�H��B{Tc��+Z>\��8H��{�\�C�#����@sX�v�:��#�I;��+Ju�!!��� ,� GodK�&�Y��ٳ~PA Z�����ĶY���Y7yD|�o�w���q�q��Ty �ݺ:��l�$�T�ԋu
˷R���TC�Rc�S�?��8�_21��S)�}����ĳ�Uc̛��+6q5o"F2�=]i��[�&������7��d�)5�Xk|D��h�ŽF'���/=�1��uA�Hl���_W�ŔY�%
�f�¡�:;s|��!sU��������l�[z#W G���fIV�փ�	�/�9/�h_g�=<P�S
|���m�b)�b�m`���-�}wE�;��V!���%r;'��>@��J�E�LX�:U8�EH����G�a�˳V�%�G�Ôh"�F�2.��Z�	e� ��ԗՓ��ߥ�퓼f����L�C:X� B����L��a��j8��&H�.x��)Q�q����؄����'��~��hI֯R���/�(]���q%�R�ί�!�t�p&*tD��[�ic ,�����`���6�w�M�̧�m� KR2C-��,�s2� ��8�{qSqF�0̒�>���\����S�1UM�c�,ӦqXv	�
]�N�T�x����s��b9��M�:aP��m�_w:�m�$�q�4t��qP{�����N�r�s@������~��������?;���_���zr��|�i��V�_F�I���O�*s�Ȅ�/����W�^�(#��^��k����*�GDl��r/SW�x�e��%��2t&�p�׳����s���D���z?\!C<U�C�e��ߞ�r��������D�!����~�Ǫ�*)M7��� 0֬�(j��i[k�߱��ıo��2�˗t�Fg.� h8�Ж,��wu5#�eX�j�0]X�34AI��%�yP�[�؂] 8��C��S\��Ψ�HH4��)_�Ğ60���
'��는�NY���4_��m����N:��D,M;���0��71�1v�=Ƕ����`p��Q@��~�C���jM���,G xߪ�;��D�e�����)v���{O~)r��-�>�,��B�/FTN��6���V������<w|,�{��>PG=N*�)�d�#�%��F<�m�F����y�YV�\�� |\�<͚���|���ER(��� �l�"��6wW���������-UU��7%���Lo��E\t���:��gɩ&�9� a�\hn(/=����B�D�p�?�]��#�����DKI�l����+�����Q?�70�Pjm9ID�	��!�0�nQu��Y��|:��,�!<�F�{i��;$W�&|����z���ڐX'4�7��� ��K��Ibl�졖Y��k�dݻ
A2@�Wz[��`���.��qM$+E��a��w渎[턇>{����zR�>ܡOUiN	��o_pl�@F��.țDܵ��?&�P}��ͤe�MKH���"�eO�M�R���?R��jO^�gc�Θp��P�¥�@�!��LHt��J&2rSB��3�_P�"�.P�h�"� �E�<���uq�IS2�A6���[m�Q��!H���8��V&"��j���c�U���������Aq�8.k��N�*�HZ���r�_�{��A��ǡ��J���4�4�3�=DY�@����-�HFBL�Mޔ�:��x�]8��B4�3~��x`؈�:Uk�ujth
�8yl��nkb��C�N�&��}����u��ԇ<-&:��~W�U���ے�I�š���e�5X}��A&�l�-�T%�_[P`��>�gա��$R�{�vV}�M�߂N����lMo6e_�"D��CH��M���|�F.��S�����Z��4���ȤP��{�/���<�:?ע��y(�h��@����!8]�t�{����]E@��/z��n�%�Ay@�2-��u�9���D�Կ�ӱ�%�}�p�=ecO��ɢ	���WM��HB�!�nY#t��w�xt��w'�	��
���4 }�ˌ�J��k��Ua�'��p>c\�4���k˱1(/�_�����faG͛�Y���4�L攎��JZ:�&��o�/�l���ҟ�#�4oo�U�3w��U���)-?�,,|7�N��#t\i�������n�I1�����88�#_HXq|w���W	86Zso����JT���hv��F҉�\8��	\AbVyȘ��!32 b*߷%v"�JiJ��[��I�^� sx���ìw�6u7i�N(R���5�[]X��V��e��]$��lw87�J\�M�PA-ء�Z��������k���۷��D_�n�Z�L�^����"��ݭ����zKӶ7����{�q��_V~/�'���ʬ�>1���$�ċ/W�,*l���^��F�Y����X��/C�	d�g��Z^?a/�=�TO%a�'�w���_0Yˇ�|�S��[��k��u���[v�%>^yḄ���U&�_�WS�@l�͋�}�,�`>�,����m�E$T������/K_��y06���X&�Xo��V���%&����E7�:���S�q����.�� ��NG�������=� I��e����w�ju 9�G"K���E�"�7%� t��3����7p3=X=������*����T����{;Sqo�[��?�y���d�c�����hp�/}�ֿ��,{0+1�ל��M*&�~]$�oaf	�vU@�3;����fi�4X����#@�/���\��P���е�|Y����0����~rC�z(tA�t���6�}�]���ֿ��QZ�Q�����
m���/S�e"q�Pb`���6Vu7X�A�pq���R�s$kY��,n�e���F,���랝�����s0�6���,	=m��T���du �[�)��+P��e��֙��ā�/o VX��-t�j�,�Y_ۋd���q��S� 4��y��B8��3�'�߼�T�l�m6p�s�e<:9c�u��b�^�eq�����D�w䪷E�Љ��,Bu�Ú�~aᅼ+�-���\k	�d�:�=QvzDI��ך�������tp�#9G��j��}�n��ZB�i��5�2#_�1~�0��r�U�~5�T���!����H�~* !�!���ãY ǎ��3峦�����*��^��T�#�A7)nÂ����Y`�������g�{4#~�iz�a-^��D:�uG�MB���~z
�G�� ��]ڰO�%�0�(��)0S��Oo]Nα��ge`(�a��+�;��&`$�+n���2�Ҧ�۹?�I'�+��$8��G�=^�B�jbߙ4��j�ݥ��T*��f	ɩ?���3Hƚ�7Tx�����*��eTS�{9'얋L��ʾ
�4�Ǫ�+(h��GUR���	�_�[��(�P��My�B�n��u��Q8����!eoR��={æ<u�m� �G�\��Up�T�(�(���-6�jUh>ʰHuL�$��
a��{B�L�Dz�X��厃��I��` 0zV���f��r��4�����\q�P.�i��,qj�?�G���E)�m^P�(d��Jc|�n���jf$��r�m;H�u��E]��f�9���\�[*���N��`��[��F��?��%H��^�*q����D��8�{�|��C1�4�e��W���g�y�qP	x"O���9Х%o^аl@��'��7��!��m���^!���淧�ɩ��Pc�0��+/x������uf
 ;�S�ۋ.ʞ:�������n8tY����Kh� ��ؚ=i��Q����w+����%�SVC߉�jM,�F��E}����H�O[׳��/�WRG����G��=џ1�,r�'�50~�C�Ὼ�0|�s����ɷ$�A[iڣ�J���!Y9Y6�~v�Q�]$ke�k��"�({5���/�!�Q��ק02S�/״�rغD���,G���`�ShێW��;��	%	�t
p�P�f6�h�p���)N��(��RH?��}��W������+$��a�����$E�n3�!Y�C��B�O��a��Ά,-RS���ѽ��K��M5
���x? �R^(_��M��j�F�婟g\���^Wh{m�U�%�EY#a��9��܌�m6�fn�}��q������%�h�|^����H~a�I)fd�ˬ�O���WN�&���P�yM�vs��%J-�{"Hg����C<�t 8T�5ֳ�K"7��E�X�ȶ��>ѧQ㓐���=��]\�ed�����Z�ٯ�v�^�4��3o�g)A=�pJ@�ok���6�<�����G�R�*@ê*�]�bM0��F��7d���~��'�eϲ�ކ�j+Yt+�8k����A+�U<`��g4��m�B��'��� �O��"��(�n4��m����!Į~- � �E~-#_O�ZO���'�������n�΄џMIG��~Xh��Za�V�v�X�"}x��%�}@��=�ѱ^��Ȳ�FI��'_���)��$1E����C���H���>�ғ�� Mß���퐆{��C��mg��t/�B��@���=�۝L!�AN�rm��F8���ep2�Zʆ��S\UL�]� s�h\B�ݸ�q�����6��[� �������ʓ(�}[zD����|"�m���Q}��/��rI�����q�)FV��;��Z(�k����/;���',_�4+l55���%����������m�YR���JLC:�((y����A,�M&-�>��I�c�N�J�c�r� E�@~{�֚������`�T
���î�~j �7�m��O��+2.t\��-�7,?C�1�l�3*�!�{,N���u'�� �c��;q"�E�{nN�=�^��vP%l��a3G�]���l/�oQ2�Y �?)s�����j+>WF�e�0m�w�ٓt�bt{����*	�@��X��_B�C��7/!�h0���r��ӵ��T͑�4t�!~t���@m�<c�>��K����󳮝�]�@E�$'�r�g[�˟Q����2�����RN��k{ۘ��K��ciX�2-��b'gݶsi�b�1Y7�@q�x�vۑ�usx8�@F���]�A��kz��9���8��V��o��|f��E���������
��������*��F��.:��Yǀ�� `�V2�XL�
3�nV�.)Jx�U�Җ��v'?/tՁhR�,Ҹ ������A
s ���]�q�ί���{e-��ZW:�dyJ�t�v���tA��Z*� x��Ț�ҧ�?�Ҵ��h�T�N���{&�7/[@�v�<�-��ƷPK���1��܊y���C	[O���VŬ��;V���G�RR�\5<�A�b�o7(���/�w��&�6g���~sƊ����S�,�[.M���{�kq����N�R�yư�mɏ��0z�>�B�wԄ�o6Ո�w5ІΑ�o#=�1〈����p���^{&�'0N�}>N����~���+w�=V�'����9���V�)�����ٰ,�	�! H���27��C�*�A*�~�1�l�ԏg-�sE���XR�����{X��u���5�f<ʹ�aTO=%ejØ@�����щ�&}&j�ID����L��e(fO��Y,�lr���tH�ӯ㝄���J����F��^��Z7+�,�MzG^�=F!SA`,������8/�-*�OП�0"�������@���	�m#į�[����q�c�YR��x��6P�m���ܭ����R�ڄ��o�ù�v��5!P�N��GQ[j]���3ڪzwVVh�&x'Y�ޝ�+���&>u��|��l���-�qI=��(B��Ήs�g���|�F��䢱� ���#�}�'&��"tS�������$�x5��g�*eA�1L�����\��R� �&n�y�O�Ό����t^��F�$��V/,������8�{��섣d��Tݜ���A6�N��<�%KW8�n"��J���Z��hY{S�UI�����3�,�!4
�K���e�X��]��Y�֭��E7z�@�q�ȹ�����[1�Q����b�����Z8�~춏��M+�![T;d9���ί�*	���w>$ڣt������쩐N���R[-v�}��lPOm.��9&:�I�O<sk�tg�M��ru�W�ǌ4a�L��e��3�6E�27����G@�t| 0f��nCw�x�v�Ӊ`�-��n��&3e����A%J4���'��g���dx��{��]��c��Ε �'�A��8޶\�Ƣ�� ������F�	}w��ϼ��RQ�t;;����Iߘꤐ�[�B��E�?�~��Z��&�I�|�V,?��7�5&���qd,��\g)�f��{z��Be�D,�\{�b���3Ȱ?Q��z���p�Q�/���_r���kFQC�Z5Zg �A���_x� )��Vwx;�&Z�=:��y�;��µ zUC]��%͈���bHdZ�#]J�V�`"0V��f���U�,Bz�K+�(��K����:`���|�����;���E��
�*���\�#Ճ!X���M��0'��d��#�"�5 � n�q�E��1��x��{�4�]Q�V�K������twYm��cZEF�/G�S2�ڒ���n`�Ց�5�5`^��g�Y1�"�C1����Pć"��uA�o/,�<� 8m�3$���H��|�9920�D��9+p�_�9����k�%4þDc��EUw���\)`\B��y���&:��~�B)Mv���ԫ$cE(��2�o�YrҺ�Ψ^3J����i����W����G��[����e~v�=a���l�.������~��e�'I��i4jT
�&wi��z����.�4����;�?tDE�4�ԩ�m,����)�������)�́�`�:���������0�`��Yz|�����n�iq����+d�sz>�W����0�:��8�oA'yg�s��`H�"s�n�拉��4�)��:���6��ίg����3��F�l
[O&��{+�W@��v�����yң��gu�Y�|5�]�f5}f	�$J����G!-a�1�fq�e��g�+��A咋u�7��T6�Z	#���Aג����F� aFP�ƫX��)�`���j��Ԇ+)\OHib~;� L8^����zʷ&�99v�#�rVl��)5��sYX�3���9V�[ǰ��W��7pb����M6NcH�ܠ
�]����ǭs����D�oR6K�tK��k�Wם%�!�LjɪQJ+����h��2Kҥ�&�h�_��%W$�8ޢb�t]M;��ك�
oT�kQ8�	�c����gcgJ@T;	C�k��w`��Ƀ?	�[&O��-)��\��!
�a���9�ϳ�W���~��Nn�7��`��gpR���vh���Gq�4��'�ȧ��A�� *f.�R.n��"㙒h&-�J@l�k,��Q���e{�hxf�j^U�~�j����#ʃ���1llH^�YG�ҭ5˟M�����}\AڦnI���^~�g6�]UD��w��ɲ�BM+Y�\���j�[O�X�W�6����R��A�݂�WA���W�Lx8����E"�kpć9��l�S ��p�3�S?OH��M�f�f��9F`c`�+\�Y,�/��Е�\��i�"�Q�����+�̄��c/�v�t�#��LOxJ����<Ԣf՘���#��J�!;-PZ�iԾ�_�^�5����y�6�tF��П�! �Pڜ㞍C$��¤7o_��/Ѻ�ֿ�&R��������/��� c[:�,&��<س���}�e�,{��/>��o�,>\wT���� ��f��2��g[���T�;�l��
 �9�S��ړZ� �ۇ9���EO�𔭑OQ��,2�4���dL3x2?����D��Z������f��r��>|Q�'KZ(�K<��dz�nי�kN�y9�.<�/PbE�5Xķ��8�j��$4)C��@n�bM�/��t�~��]O"E�}V��Qlf*w�YFI{;�ӿ�M^ɷ�S�2�'0�&�k�R��1�zlcB(+ 7�5�e��N*+�gh�=c�c�P�6"bH�W��V��I�	�/������q�NW���$m�M:<B̬��b: �(�;hM�QgwVQ�GB�W��!����5��)�ҧf�s�;)�2�Xe�d�	�>*D-8�ڻ��O2�F��Ep��#��[ޏr3���@�Q+*��deӃ�֭�͒�yN�_r�zzVl�,�t& 
�X�yM�I�C@1�S#��sK��ʉMH�@��HM����1D�ew��
soQ��7�d�ּSm6Z����G)����<9\���p����Hy�@𲣐��.�A��/���J��_�_��|ُ.�TZT�� U�Ú�o��ȃm�v�\���5y�^�(N�i������=���׵��K�Fe�7��^�?%���}�ٙ� T1�.mW�o��[��ݍ>%���+9@��$���&W�l��	�Z�ޜz���"p�?NݕW�_&�Pp��0�4�y�MG����|ϢX,��
^h���&(���j7X��S�E��(͗s��pxY?M�������Ǵ-��0�=�Kb�l�?R4%�<6��\�j걋����/�We�����"�c��bo�͞gA�aú,���Ҏ %��D歴�gf�*���>�iB%J`^���DQA9OO_������x�u+M�۰s6?�F��B���
��&C nqYN��2�R:�4g�z�|�a?/��-߳�t���Ȑ$m��ggIT�^<� �jly�H(�hX9���T���S�y����_ؕ�(�4+�)��Lc2��iD��!��'�($�i:�� ^N�vGyz)����T��,���0�d\���G~�$�+/E*�����bf$ALX4
�{�5~�5v�qM��&��Q�_�WزGj6���o���S@�ta)��i��y:��skߓ=��~^wh�VK�+��z^��Ơ��ɔ���~���# 1O���G���ޤ��XAE�#­2���[/��۸�w☝�z�gH\�R4�+�n7� �B�����	U6��2
��'��~P.C�೻������iC����Vr3��3v��f*_$%���a��蠵a�Ί����oR���T2��;O�����~G�b�����A1	�*�
���+���r6�<H�F������OB|1��Qɐ�l�ƗkP��Sv3���ݭ�)�.��P$;����K�B .pv��]�/�!z+(J�)ޤ%_������w6m��B)�D�( �:��u�/�l�������S�K'����0b�jG�9%m�����5Z�L���'�Q�B�� �HK����	+�\����y�{u��b�a���2�yXmzЃ������U8T�É$-���#J�����ϻ�D�P������剳�^��������D!߾�2�����0T&�㵂��a�,��g�6zn�py�TQ��q�i�5����o���1��M8�ȕbH�UΩ�C_�AݏK�JA�� ]¸w�z,���ȝ?5:����c��g��L��,���������� ?��w���(+MU��4��S����P�!���p�
4;Vv�ű(��	��A]��~�'.�1\������9�oEUԳ�?�
 �SE�!��l(�gPt	���V��@���t���!<�3�]���ЄÂ�f�mѹ��7�
�?��;p�G���A�}�ANl�푥�����]�7X?$r�ݯ�}�( ��Y~���1�X�6�a/j0�p�����.�Fs�>j����&姲�dx�+Q��s��r��<�_���Uk�S|��i^����<l��?P��콤��U�Uf! +N{��Oͱe+��ϓm�u�� ��Kyd��E��_h�)��U��vh ݫ������3�m��S�/��WX�,��'��F�\�~:Hɵ�+�� ��>s�Xu�w΍�|�}@C��R��>2�)��(/�9A���}��蘉���ʞc��Mj0��+`Uk�'��[������-������PݒӐ���l�L�%��m����H\+�$o3L�&J1	VbP��H�F�	0��zte�|x�fg�u`b�v��O��������E�T���z]c%I�T��.��X��RI�Qc�ʖ�p9�P����u���e��:Ќ�`m��BhVf}�&��D��&����EJ�:�S.����a��3�GȈ۲�oՐs-�]�|��E��
h0����i^�K�+k�Ics��MJ �Z��	�3�+6O�S5	���wʙ�jd�*�Bl����9�<s�S?�t67L}����ڣ����x�L��.dz�Vr��_�l��� ��Һ����.5�0a+�����>�{aq,�Z���\u�ԥ���dt��!�1�ET/�ӭ�������K�;+zɷ�`�@�QQ��M�o����2l������d��7� t)j;Lf����F�)Y/�]`PЮ?�/�l�#�O�`��b�p{�x��N�?�9s�P�+/�MA��^H�������!M���By��� �$�/�Q���Pa' ���V!Ħ䇅��)
���lMJ��F�h�0�aas�]�����:�&��B���^IM@��^>��"�(J@W>Z^��$�:�)���7�GU�������[� E��w6>ڼ9eaȘ7$�~��.Jȸ_��[��Z��%d�f�QhT�$%9�d&c����޿���fx�q@7��r���$S�`�
�QT��W2��}�@Ԣ�;s���1A�*��2��.ɟF��s���6�Ќ{(��e���x��b����p_� ���^.W�k�sjm!H�-&v�g��}�Nw�W� �~�X�j]hJW�Bʮ�Z������������W�����(I.U�u�lR�=q _�M!���b
�HmN8���2�%U�BRC�-(�n��>�3�m�J����`+�K�n�����H�Vq<�M�^���2�W;�.Az6ֲ�L(���J6l��([f���jqem�6c�vQZ��he$_�D�y�D@ʎ�����\r:;��P�$緁�`��� p�����<�9�>f%׀�E$irud{�E����&о:Y+�D��O��=6;sk�?T[�	q�J߂ߩ�]�DP�# l]�;R�`(�R]�w�7���	ދ�9��`;aH4|�U���i�a�f] -�wp����7�]��*.��C�yC�����f�I$q*4�?h�I&zu��Y�ʇ ��L�ױڤ�ak��_-����8]ԯ�2�CT�U?,e��׌H�?{�mK+
Y_Z��me�Z�07�q2�:��:�D'��Z�^FO� 5�����2=z�'�U\d��<j"�.��ŗa���9O��}�'7>j�{�!�a�+���Qa����B����ez��� ���y��IǞ�8�p7�z0�%L@�1�����	Vd�_D��9JP�S���,ϩ�|Be@��@��m��;�ek�O�]�WM跔���@�˩x`�[S�t�U��;�u��׈zk3X�dE�]�/�?h�e�X������sq*��V�ǜֱ��3[����g|���+���M6Nb��#Z�)4S�Uv!�`u��B#�ݜ,���Fc�K{���=�fP�R�����4�f��7�
�ya�fm�y��VZ�N[V� &� u�NC��r��D����{��ĳ7�B~�iGu�}�ekDP9���t��T�o��Ռl�<�Ǹ��dIZ�8���2����Kl�w05��&�bT#����oU�b�A�0'���!(tQ<hL$����A���{*�M^�� `����K��^o䜄R���\�+�d��r�Hg�(�]��,��0��?�\�1��+	B�Ǹ��I�^���un�P3��p:"k(p]�#B_�?J�s���4.&G�1^���f�rٴ'� !Ջ��߿x�p�b~\�Nm��=y��w�*� ɼ�k�$����$���y�'���dм��M�A��W�eb��h�4���f����
<��q�~���ý}0>�4��z"u;z�>��wf��qu���@�Ȏ����n<�n��|������eZ����)�
�U����י�*	�����9/Q�-����_�%�Ba���Rw���m��J���0k��bo��[��*���
����A����c��d"������,F����M���w�M��n�����yfS��"��*�>���	����I�x	�׼���o��q�]��P��'L<SO���xs����f�d�i7���L�%;T�ym��}}�cU��Bv��AƿXG�ܣL��FI���
2Mڌ���Gߚ���������:�ٜ�w��S�����G4ܜ�]b���4��� H�y�et��Ok��*	�K~5���Qs<y��*�V[X��G{���H�fS7)��x�jQ�k�6~�`_���,y�sϘ�-J5�dTG��:u�����n����^z1��ڨM��dO��C]+�e(:߅�bD�0��Mm����ٸW�D|�'bmM����V�0y�!��2�A.���P\$���R���ӑ=?[��v�����XC������h���eSsTQ� �Jp�^t�p"b��.4��\7���j�g�_y����`3��)�p�R���)K�T����������Nb2j���0�n�z���%}_s�vh���/l����x=��'>��g}F�U^)��V�@���~�;�� l���u)�5#9����"��eM�*q�:S	��g(���vW�C��+�C	��L:I�A%�.�g$�Yz6�vW�"�@XA�y@lfE�<���QQ���[?��T���g`����="ߛ+�.8o�+�kv�1$tsN�<渥$��I�����g�ٵ��V�Z ��@�[0�[��X�����-DO9'�)�(��
.`9&/�zv�<���U�%�p)��G�pwYp���N�'!�
*j�2���m�!M���9ԓ���帣$F�����~�B��Iؤ�ĕT�7�����i0t��'�;O ���{زe�p��>=j�Z�Js�������w��A#S�^w@���Ն���>�5�ŭ�7Ɉ��^M�ӂ*�e
Xf���e������)t�	��КY�a�C՞޻;s~��&gP@�A'�w�vl�����2�!l����cY�;�0�n��C#f (�id�Z��q��5���A��	�Z�z�:)��\�).���XOh�,�F�)�;F�	���F�.�(����XZ�2�!�����o�'M�{*����_�t����]&o.,��zvB/��GHq����x�B��(�YZv�YSƈ^�Z����8���n�5�D�B�1	"���86(G��ڣ���X���1�5Ļ���pK �H�񥅆�ge۴��k�]��f��R'���q��Nm��k��/�2��@�x�`҅�t�U]�ЎZ��>3�j�~4��M���1�u�a��{>x?�}�1�����\�����3BՒ.�Q�{�O{��Zr�(�v����i@KΥ/��rY*�������z�p���F���1�r��T������%\��W�9�B9eT������f� <�(���ɰ��^�uW��	��}���<!�$|�2u�x������$�~Ҥ�%�X�'D<���Nd�&�;����E�	h8��%���O���
d�VNw׶.��4�{��6�íC=�Ä��"�E������.�Q<��r]���)��^bk��RHfR�I�'8k��BIv��"��I�Sx�aLou_T[�@�)��g`�KwD6�P�V����f��Z.V��|Y�g��|tx����*"��%�>8J���̟�5	��A�����D�gN눨��7�>��1������L"���q���Ǘ�Y�N��8�x���������.�;7��b����Ʀ:-�,q�A��-��;��7(��eϠէ&�Ի��Cf��o�� �Š�EWT�z�R8_5O�? �����	:j#>W�mS�8�+��i�ݹ&���P�[.����,�d���o�W���\Um1�8+ٳ�fHӪ<*�v�G蹛�F$и�?��k�|�y�z�ZɚD�MͱFJA�-���VyKjhĘF��#�1�@�� ǷN�6���<�u��^��'�Vw�O���FJ���7q �|����=���u֐��u�qÅ�Le�"h'm�����Q��_�z�N�?�f쎆��-Z�9z|R���qY�R9�ZR�I�y�J�'
#��*�BS|t\�bpf{qb�kC�g�*ÿ��;CMpv,�͜^o�/�a�z�Q��5Q[�=��,�de�'~�����h�iV���v�'��[*Ϻ	� �fPMx K�ݥe��@^�!����5�����%��q�XBSpI�8�����3m(~�ꚰ8��
+�u�o��k��s��y�������su(�~^p�bi鷷e����6��P��7��>��&�Q����hA1�̻�RS����`��u�$(�[i�����]��C����M*n�G�p�/d�+=��'\��8�����i������V�)�g���8K�mqX�w��+�|��*��$ϻ7��rC�Y=f#�f�<�5C6K�kRΟ}��/L��H��8�f��s7
�������W�I�ܔ5��&H���Y�*~q���� ����	�6[=m~�L�.I���l�
�Y}�+ѹ�|? rh|��{��f������J/�\��>�d���<KNy7�v�������ߪ�?�5�vYH��~�\6����E�ܳg|�e�r�p�{�i��pu���qȽ����e&�6�s�x���;y�S/��՛0��[b���Hz�i��W�d#�����0ŵx�NЖ��ٷ*���E�&SWh�!N��� �2��
����
�V�+�̿�<��O2vK&�#sE���-NӲ�~�dbB��QU��]�m޺������hZL�1Uv��2F�;<���nh�u��++��ັ1�#�����t�&��H�oI��1]�ʱ�9Q�=��j�����~�>�tg�_!��4�̆I�h}_��Fm.���W���'3#� P���G70_��
��.��Y����~���(RL��"(������ţŌ���G�S-1�JJ�b��(v��٣��ӆ�f-��
�v�<��寺m����6a�U�U)x��m\��EP(>���E����� `�V�>xvK�����<�?XN�E;:�!��!�L���}�H���f~�U�Hmtٳ3�e��!��s.�yɳ����VU	E�;~�s�|uq��2�������V��S�?'V�"-X�E��{�pН�AX������+Ԭ���c�v[��G&߶���@�o��
n���2��OϏ�����V�����%��hq�R�N���"Wn Z5U���7v��_�9#B��If�z�ϙ�*�'�êa��{���:^C��Q�ZmT�ߌ�����[��t�e�"��n�Ç�d3��
+�amzj2�/)���r0�] ����x��E\{\���3jf(��<6�h���U�.�����'�iN�����}��w!N��H������V��<�Ź��(_!������O����Us�~��#g4���������f�j�z��:�	��@yg��:��e�V�����x�G�S�v�&���GW�-U�u�n�4<>0Mo��*��1���� ��*�m>�I� u3�F�X���<vu�|Y^���8?筡���%-A�0�����t>)�� �.�����[]��/y�}���՝��nrp�}�+�`+U�{�wI��k��N��c&/�b}4=���r@���J�6��w�����S�f\Hi����p7�_@t�JE6��uYLO��)j�fu�
���Ҭ�n*�ѥ#ur�� "5�WIA�#>º
r���2B�b�@�Χ�T\�MK���3U�e�4�����n�6��W#�L��	��>�3/�Q�5��
����^�9�F]B���o����B��l�{ĕ�"	��z�zY
pܖ�ND��y(�p>ơfU����"̱<UMH�oY&��1�7xI]E���� Im���6�)xǉ6ѼNcHl�`=w�h�fٍ�ۚ���	�m�S����7��Y�Y�wD��~QM�և����b)
�3D�#c��]d�܂����"؏��P%��H�#�
v�"ʖr����� �6���]��ء0�����(��'@@����E�RG��╯�"X�ad����*�#
�y��/u�D��mM�Qs�sb�0�2}w�O�� e�8�v3[�ذ��X�vg�h5�S��w]s��m7��$8rŞ����k�}�;
7��C�e�v\9 ��{�oaW��#s���\F@�Zx<�>�敡B��`<���M�T��T�"[HJ��,��<�,�zx�3���\��\(��1�j�y�%�W�N6x�q��"�=Z�݆I�Q0"�3��3��0o�
�����n#);y�P��pi��>�vQ8X.4�1��n��H�O��2��	�n ��W���ߕ��s���c��mwi��N?d_$�q?n-�c�l�e-��~�$�\��Q��7.����@��S�%1ȹ�<S��!���Ǒ�{gRdl"w�l3�ǌ�M�{�7I��k�S�2�z���>��_f$�R#���3�+� 9����)lQЉ�jÏH�,� ����C��-��6ev���r�̭��arp���tH,bU�z�����~~exe�z�v�P ����,�<��?1����+�y�k� zI�%�T�����*�������M��鈇��?� |��ѿ��؋����q}��^H�΂oF<�G�9��"�9M,��h��+WB��ڋ����/k��%��֖2�2�å��G��d�?�4R��c�s�֮��$SLt�>8�0���:��?���s��-�|d���r��D�`��*[������Ջ�v�+i�7�`Ы���ã/�FG-�ψkޅU��H��<�ke�I{�Dn�`d:<�h��%��Z��=>j��Ɂ[U��dE2��i���������}HmaJ�k��̖>:����Ԍ���z�OJ��z^�%i�$�v�IL!���s S�Rf���}W��0\���8�+w�gO ��T�Kr:�L�Mq��_'�k�u�K�`|n� ���ق������n��ڣ4r*D ��W��iY2��Z��|k���;�QTw@2�n LX�QWK,�1�u�\@�)!$���ϡ�kV���N��YԠcԶ����&�;;��x���"�7zyS�^��qTv9{%� >NW�w�0�{��[f�mZ��(zkz���*�z���} 'Q^����A�!��W���8b��"�A=�NB���[��a�o_c-g�K!^3 �<~vP��"�A�Z�^K�ᳫi��a��őټ����7����W� �eb&SR�����H�Z��5bhLOv=x	����Hn��X�`K�N@�����ʝAo@Cjb�f��}A�)E:��Ɇ-�g���W���]m�u�z�ׂNN}�:\�l���td�{o�u���?��5�-����,��n��+����S�)��[\�̩w�J�:~�%$*���:����=�^�Ը1&�Ms!�紫"�����rjL>ĺ
���;��?&
��(p�D�X����EE��ZUsA��A�6
�u�u5r�-Ƙ`��!��v&��Ng�C1C:��\��P��
��e�+^�{%zT���������.u�Nn�7����D�zu�O��e����9��7�?Bt.ϥ$_��&w
��ӌ��{�3<+�����+H��jBCO��e:ꅆa,Ǒ!��{��G����q��N�?ѥ�S�e����n��W&���F����k1s�AT�����L�X�%�/��_�tPA�%�5t8:��u�hq�q�e9%��"&7.<�s$��{��?H~��)�4���mc���5
F���̫�<?�+�5�N붽[c�6�{Z���>y��\D�B���^��J pƟ5�"�a�3�n�����ģ��2�!E`��&�*��B����O&��?>.�zD�y�}#795�vl�
�וY�*_��ys2���7�Y������	�?2X�d5��X����]Pdz Ũ�C���ax|Jz��֑�jh��]�-K�-����h���I�"��u���)��Y_�	�S;G��[��ա�p`fTR@I-�ƿ�6[w��$����)��6D*Od��j�D�ս�*��䮌|܂ow:6��ϱ�{I�����.�%���C���u�_`��i������=A/��]�o�YĲ���k�Ѥ;H���q��%�!�(�H�/�ic�1oYޭ�pO�탸D%�AX֭ݓ�U��U0�z��r�T(�ov�XڊW#ב�qf&ɣ*I(�"ST4�%�����t�a�^�:{-�*Ëv*��p>�ʠ=���^Un�ߺX�%&������[` �z,쐾���[_n$g?US~�-,y�����8S$��"R�.�����m�4Pً!�kӨ<<@�w�r�|"5iﬦ1��x�:��[p!0�ҏ�{"��^ٰ����T��ֹ���o��!u���Л��y�=?��u�����H���E= rf�#��̥���1'��NI���Q��i�2J�=Lų���#�D0�ݟ�!(��u�*�B*Ӎڰ���VrY~qC\���F��w�Lx��C.�����>d�M�O����$jtң�9D�jW�ԉ@jIA�}�
����DI�(AAr>,�����G�cg�#��Q�!��:�T���f��h��[�O~��* )\jD���C�� �<���xJ_���bP�AQY� K�%1���iW� ���Mn�Fڒ�_��@�(��*������������P#�(�,�7?�1�?2I�HOa�mEs��<�?R;�V{�� Ck���;�#�5�@$�]�q����U-�N�#�*�y慎�R���a����-�.��J4�En7�_�o�N��ɪ�����C�M�N���XET/�6��k� ���ڍ����S�ز��ߓ�yݙw�Zx%R6�&~Bފn�M�B�%r̄TFo�5���2>���T,�IQ�At�Ȃ��r$�*�{��c��fL������ڮi|���c_��=Q�6|�֠�'�ۜ��T
_��R��a���/#�'���_a�0�1��_~>'��v-�$�;xAu|O�]�g��
��XhS����C�[�Sd2���x
7����9�&���,�@�=+���=��MG��.���0	��a}6G���c�	l�'��D������Y��	��Z�FX�z����g�®Ù�'�X�x~� ��$yz���c�I�^�ı�T��=ۼ��&Sh��Fr����rD��n�a��L�}����m�d޲�;~[T�\�΋�iЏ���l���A=�R�:��k5��zu���-�kt$��9��G���n,�ۀF)ZŦ��m�QK�GgS5�&�h���/�]���.�{8�W������ `�y�i��	��uO� ���0�2����]^�sެ�j�,��b�g���vw��h�V�]�6q%�:�N@��-�a���/�U:��*��� j��R܄�t<�j��Ԁ��2hā�:~��e��6+��wc0���ٕ �cp� �4H)I*mXD����+J�̮
���޲��@��U+Ǭve���>I�#����`�ؼF��~�	wy���^�UD�����'��z�

_,m ��{��� ���%ֈ ˖��ߢ�*R�6U��h��'�Pᱍ�{V9�΅�eb����XP���6~H���;	λG����H��mC�82���3 #-8���#�=nB��=
��3z��1Q62Q�B. ��=H��3�=�0×z-��0T@0�5=��Z+��r>�`ū`=���P� �O��������0��Iwh(B^��B9�BoIq9��*p2ü3P��؈X��(?4=X@I�����e�&���.�Qɮ���3i*�|@�XJ'��M�vn��c����t�Om�Z���w����I�+JF��a��Z|}\r�����v?��j:Cc�լކ������*Jfޙ�/ԅX�oK�q���f��25L�Z�c�/a����y����f&Y���Y���e�K���Bep��'�����&Ie��Kb�s��'�yp��1BO7�C�~���H�f�B?)q���u� �@��x�� n!�]h�غ28M>���!~�;�N\gh�����=r�M�G�=k���L�����>�hQ��5|A�5��$��[��G*T_�G8�� .��	���H��K7X��������9"��CK��gd�;"��Z�n�Bm͗�To��Xu���U��y~���NJ��8R��!Y|���������	\`�v_��\����6���_�[�zJd�L�4z��S(R]V�~TӀ1�ר��/�;��?�߷�َ��O��]�k�4e5�%]��u�sؑ�1ӿ���d�r�<a�]�kM=�PDa��o?�Od��"� X=���]yJ�ad�+�:!�]��_Z�=�`��] u�**A�?� ��dN�3�i���A�c�X�A*�k|G^�j|Deτ��%f���m�V�}]��b^���Ma�G�,;�5�w�1wN#T���UF�q~Va@����PRZ_F�Ƚ�O�ב)�^�=ʞ�eQt�7{��y�A�ݰ��E���y��~���ߝp������A��T�"�$�2�9(�����6�v~A��6�O�7�����Vl)a�Ȓ������_�ޠ�lT���̽�ܭ�<
|>Y.�>�h� �h�x�pm�@�U5c�a�H�ꬠ���ڛp�֤��(���W{�1�jcN��f�ۤG��]���&����W���U�b�%�(ө̄2x��L�G�x��Ĝ2fk� �q���$��~�sg�9$3�a�"�*EB��Z�fY�@����ܓ3>�]̗��n|�n�'rU��yzz%��)��S9��;eBE�YS �]�E;,��8&u�{;���W���*d�[���(?�z��&���'X�V'��Ƈ-��R}υ�I�	^P739'����ci[G��߃���*�Sv�槯wkjÁ��$i-Bǻ,˩�=ap96�Jl:�.4 �i��I�'��ij4������Z�ᥦ2��~|��)eu���PЄ���_(n���/�ڕ��L�R��|gw���5��ƞ#��s�B˞���x���l����˄�	��B�t�s�����)ҳ�z�(�4�Ni.D�*#BL���k�cŷ��ϡ�&u��5�C2��8�k��G��a�2���(E��"kB�y}�&Qt��k�QR�0BO�ʢ�W��.e��,�������\�_#�G��mM����2���9�������e~�w�[����T�N�ʁ��q �F�V�;o͆���r�=|* ���ʥ�ߍ{9�k���N��od�#G�z:��C9X���9���8p)V'��Ck��I��o���w��5I䄛��3!ɸ�ʸ�0�T�q��C�]�pb{�����o���$^�����!�Ӷ>Vh��ݽ��7��Mhq�?� �3'M�t��a�VdʤUM�қ�ζ���D����|BcU��7���Βd`j���M���������)��
]͗�q����!5��W�{82ދ_y��RUI�����/�MPwo���i3N��j"�؜���ћ�-B�t��Φs'Ҵ�hNm�.Ro���e,6�Q�S��JxHG��S���VOg{P�	H��	j�3�!&*��ﳸF�0���n��_��ӵ�8��W	L
�q9����$�����%��H��A�i_���=l�j��ފ.�4�t2��`;�vT��\��T�"�Q8��]���l��d�P��yU��R����~���[�Z�z(Cf�8� ����l{0BJt�=������:���:
�Y��K��A���Jw�ji,�@�S�q�ɯ	��=�u���| }�M�yu����;ѥ��l#5z^@����͗�2!c+�4ǻ]�����& Wy�ߍ�L�������qj��4�^�#�"�nZPw�|���QA�s�y+6k[�J��6Z��Ƽ�p7ODZn�ya���+|�Vp��Bp�♲�O�f���fP��b )�s$u�:���w���B�wEΙ4�����Zr�#ΐ�N����	��n��J9-h�f���2����m=�����e���A�dw*U���M�[�c|¸nѳt�2˦���[�F,1wh���ϗ_�*��)l�qq��,A��q�8�� �~^jOdaNg0���Pj�V��jޫ�;}�[�ڵ�N��,H��*5����	�eY:)��~V�������)����i��.KY�#�a�й����;���uɜo��J�nrlqC!�i��������M]�fu���TuIdtv���m	(.ui��ʰ�z/���҉����šz�����)f���#���;�e6P�� -N�B����[�i7M��Ƽ	4H�\#�:.��8U������'!��nСϊ����RPH�����!��4ʐ�#�t�d5��<�� V��(��Ү�dC��A?�d!g��`c�072H�Y,䩙y���9�8�ok5�����5����cv%D��nN]}ń˲�䵋�m��ӕk�σ�����Ҙ����³�&�H��ٶ�ݛ['��0�´~�.\u��_��T���3�z��%~��(O�~�d}�39�y��e�%��K���;�e�q��3"K2��T� Ո/��^�&�KM疥)��Z�7�)ȏ�Og�d'xv���7|	�t{CdsM=�x�IlL$)��{<��]	w��$�̓��v����B���#� ��������~~�1f��ۗ"�]��]4�%�'8<$jS���������$i�S���`�_ ��"�0}�ky:;>���k�阊�6*H]"0����;�J���@\e_V�(0MZ��}�<�/��B2���_���Ԉ�pA�u��ouE�X)�s��m�JU=��͕j�B�(&~
zI����s\�X5wK��u�( �ib���'��)�s�oǳ&�綳�L:3�{4e0n���G��F-��gx<�BQ9a/`����H AUH�SC��������ɽ돲����q�B�bI8��-~��)%]\0�1]��2��/�����J�=��O�_�O4��;i��J��ߟY:!��22����0�_-�8AvP;Y��3 ��'���Pk�� ��"��S��^��f{��!B��\7ʙ��J�M�HL��ә���(5Mk�]��b�u�o�� ��HUGΘ��tৄ��k'y�'�~��U�ս-л���6i�h�C@���̀>�Rx���u(���n��.��1_�ޖ�K�ޱjD�@�� �@���A�7��6�4S�_i�ϱP=���ڪ�_ղ��r�y\��r=pR�3a��D��	��t	���j�K�/ �:��H�t:�&Z&��E�H�]-���D+�sH�[�HQhg֪ؑC�����Y�U�Y�k(���#�|����.�З�u��k��Cԉv�פB�Sz�%��$t��r�r|���ή�z儴xR���s�{QU�p�J���ۜ�U� �w�������z%��W���>7�m�˷�Ѕݚ�U�ɗ�Ń{��Ը�+5��;L�nS��p��WX�z���4?au+HvY����̣6�-j��9I߷���-�7�s�G2�`��ML�x��ʟ����~ڍ�������C $�e���ɏc��ɖι�sЊ��M���@�ٻ�&�X0�8 E� ��l���Z��R�}�
<�j���D�c��Ss�<�y�<l9�/g�g�1�Y�Uѫ�i�Ӷ���y� 1RS��!N(�\�r}��I���"�~`��g?���Z7�JIi��?Ӗw[�� �N�j���Q▅zuTP��
�R���!l�T��pރO��f�y��N�5w�|9b�ؤe0�I_�p"E��ĵ¿~�'�%bE>��8=����&KZ[� ����	{��t 9_�/�la@yC�h4^�Qs��\��A
f�Y<�f5y g؍�ը61�o
닯�z�Τ4�|��=��A�8�	C�|ɳ�=�h�!�^��	{c����S6�~���T�|E�
i�S�����#D��T*�I�w�����뮟^,�V����j�xU-Lֽ,�Ѽ/9UK�/�@�7���Q?��=�����EK�P��O�,��h���9�g�O8Ҽ�1H����_�#H�?� w'.Tl�rS����	"�8$�����5,N���a l:Gm��pu9����0�I�5[�Mv��Gb�1I N:�s��n�.��\Db�Jp e�]��G�?%��!��R�2&�؁ϭ�8c�F�G�rah���)�!1������4���q��ȸ�w
j�6��M$^�I��N��<]��@���N2Zx�&1�� �X�4<���R�$�ַ��-73x��J���r��׶^x2Nm�kn;
�~#� �)����!Z.I��
���'�d>��,�e�6�_e�2��1���ĈBN���<��i("��Ė��gu�����R"�S(�5�X�6!Jg��C�����ƳcH�I��4,<~��[�H�8�ɾ��%V* mui�7��U�����E�^�rW��>�	�Y���>���]���lR��'�*�"Mn�8�a���;�Q�ßZ�zD���ɴQ�Y�:�Ƈ���c�ϢrW"{[[~1���5Q,��܇��"z�S��??����%i!Cb�i���9��񤏀#-D�U�����-�/Nܮ^�M��#����_r2��[@,�F>�0���}���16�j뽗ۦ�/ާ7F�'�����w��<ȁo���I������k	�!�㇋m��τ2���l��<M:����¡c�7=�!�uG�Q�t�i���AԔ���[|�+>����4'z���]�yܟ+{�n|P&W��ois����>�ڀid8H�n�940�)��M�"�g��)�5Ò�Hp�t=�
A�i/�����
gKz�}�r��eh�/c�������/�hS}s̿klO��U�0s��,��/�V�15>1{���Ȉ�� � 1.��p��ߙ!A�\���^]8����a(&��=SQ���n�ѱ�7�����U�|VF�Bxvi`��;z�Z'�6�Y�V4Fin��`"!�P�L7\E�O�y�e�|$�'@z60U '�6@�S"=V�%��5� b�qE���k��m�f�6��Oo�t����@�L��V�_A��,����3�R;ɑ���|j���x=d���[h���h�l5ƞE�	)�!	��OK~��o�
ɫ�$D3�K���􈧍w��l�8��|<RU��'�1��mb��LC�n�U⤠��{����F}aGV��6����(�[��l�5֍�9Iը����c_zoA���D�ؑ����M�q�S���r�%�ڠ��H/(���D����0E�M��φ���-�3�p_�.���`ۓ!�
���_�Nuv�ȁ4��B��ݖ�Q�ʝL�����;�5�Od�`t��|�ʊy4�~^����:<��.��HTR��J�%�5g*�v�7����v��k��d��4�7��-f�d�U�Pa<�u��~�3B]����FCtAr_e�Z�X7�#ӑ�BY��oH�t"�H&I�y��Ck7dU���Q1㦡٥�_>�Le�a�_�� <��"��FmT�b�V�#�����#�a�)���ۊ(2K�6'+�rT�!ۉ�gZ	����"qo{'1Ԛ� \1�K�!Dr��?��[��s�Bp*烝�5����_�kGe%Ӛ[>Ԙ ��Y�A.${��=~�h��)�K>K�����t�#�����N�E@Ϋ��_�X��ʙ�������ߐJ�b���Sc {(�S-��,`�Lg�b��,���>V��[
�D����ARɄvF�:��w��I�I#D�A�a�ϘSu�%�f���SW���;Ր�9�Do�6ҳ1�%���R��+e|¥Ɉ�1�M��G��'OXWx�
E�D��$�s��Ѳ��#�W��G,瑲
WwG؊<K
n���3����'[{=�e ��,�;j��Du���ΠI��ʍ�9{쿚�Q��T`݅V/�z���VPo��Ǫ��*��f8�8B'E�!�R�:�^���)l*�����)�y�/T�d�'�����r G�`\Y۪����
#��b$�/o:J^Ք;��iVG�yP�Cs쾺OwD��f5=,쁧�Ŧh\��X��".)]�௒d�ov겮m�S���s��5tE�;͞��rX�W�1��	������M|�,I��Z7��9p���C	Z[A��`��ھ�x&b�FL�`��� �8��%�&:�f�/�lO7�{$/p�^��I�8j�Q��U�۱9F��_n3QD �إ��� ��szm
�s�4�y�ɛ��h�~;�d����!��q�te�*��UA6wYq�^z���^�L$pmN�k��;������x��>�Aa�MH{;��s#�CI�)���c�:+"z�QM�����hgcH/�먤������9s��t�0��,��|E�cO���X�UG-�#ʀD��xi(������tZE^+�xc3�bvV���r�Lci�m<�t���ި��䯠n�kу�M���H@J��9���oY��:x�:�����ð)���
=�+�~*
�iz�!��×�Z���0���;D`��v�P`D�<�ǈ����-�"�S�{��j�F���VY���3��f9�>������������%{�X�1p��(C�R�	B��LK� �M�p([?�l�DdʢM����z�H!�qH�;(!�D�L�,�SI�c�"de���C���Gf��Ѣ�tu��5O�8&@cx'W�YPM����O�"*�r���q������y"���t�B��\�����hQ��ʌ�\D��̊=��qVbL���h��Z�4��O��!�	E�ؿ���	q���С�-H,X8�MK�Aۚ��[�M��/?n���ڝ�-���D�xu���p��C7�N9��[��{�d\����i�$w�g1�A���8��8A�}���1\H�g�W�I^X8k"�{����)�/dy$Y[�(:�НT��I<��������~�`=l]�LR����t5ݿ�к��6��+ɆYǲlzH)3���m����P�5}��r�B�� EAf��.nzg��ix���RY��?z�y'(�)@�v��n�w� ��ؑ��!�h�0�p1鋠΅']S��0�c_�1*��LX�w���3��~d�G���%�nޓ$����F���|���7F"p��˟�_�1/ү*Or��3 ��҈�EN�p�mڐ}7�]��;�r��{�;dCnO�0�U|��4yR�c���Է����4n�P>�[�ǐ��[J
ghc��~!���c�5��1�ɯZ�SHs ��[�&@�	�~���lv���T�O��vE}�K���j����V��efC"C�c�;��ma����ck�f�
?t|�)�j��������cc���I�u"���� zf���r@��'�1�$qle��ͦ��������>����n�*�@�'U^?���L�j�_�m�E�9Ӣ��7�M��\lz��_蘂=���9�������p�������ˬ�}�Z�W�r�֋�︺Wa�[/��I����ڣ�U�z�Y�kQ�-CNX�a����򕉽�K�y������@����w���І�#�u;⽺�}#�kw����Y�/����tΗm�,�I�y���]n���(�F��gw2�_���֤u�0�e�B�������k �2ƙ���U��՛�=�&�07NT�Y{.j����#�O�I��/o5p��\O�v�O�1ݼ�	�+%��2xD7�Ü�����cy`��K�#ף3��|�"��S�VWev/rR��+J�����d/k�������&��op�]<�Y�ߣ�?ύ����_����KJ�*@��w�b��/�<�~'���V��0	�O���T�	��TT�����`F�D>$ڬ�%��#ˠ��?�����G@����e�a��?2kgӲG�F�r��o�%]�o�v��8���{h�X��ꏿ��Um�n/�*>��F�d5�P'D�ӛ�.�"��A�*�)�R��$�>���K*XS �ya�f�^$�+~ }�W�10�	$:5)����=.��d*I&F,��+lb��:�5�e��NEg��<�J��r��.��J�2���:j
<�4���@o�7?Ly9H��(y�<|����ۜVu��T�"�좟�[�4�]�]��vaS�yzY�B���.a#] �Gy�^�4}�y�e1b�2��_	'� i1/-�3��$�X8(@y��;�9�9f4��X��u��c�"��"���dZ�$E�c8]�@	�w\�aЏק n�>�Y����i&����&x�����C{,.���$�/�f3͟I9}>�\�~b8!c<�����Nʞվxj�I����O���S��S�e���n�/��<���'s�gS�vUM�'���+�D��g?T)G^$� Õ�mZy;����>|�z�_��|}hf+^<!��1�@"II����"��GD�~!�O��z��j�,� �K��������3�N1���a�Y6������q�����{��F:�V�_CUi�g����8����0�M��G&@�V5~^]])�@�.\�/UiES�)��x�i9��´�l��Ϋ�\`�3fۜo������(:�D����1���idC����=���RcC�j�#ُ��Z��O�@ܼ
���/i0`kAh��˷G0�}@CgwbT�۟SG)p�&�vk���"�����Lr��,�;	)�z8�@�1�8B�Qr������ov�6�9�2(�Y<���=�T@K�3	����3E-N[<	q�++ҡ&�5��x�4Q&���]��W�t���E+]o����N{���ݐ�ԃ��k"k�˙J�y�"w�B��\��x5����nZ1\}K>��s��I�]H-O�)=��1z�X:���f��Yh�Ue�Y����B}6��m�y��q��R��O�uT@1J�DutU+������}��c�6��E~@�J��`�Ȱ�RZ
LG8��6�eV_�Ƒ�hGT@" ���F���a9�%�Q�i�Ĳ)�;� rB�c��,�<�,}�zY``K��8Z.�:��#�ڼ���,?��H��zA��G�U�GZ���2~LH�ܤ	��%ks��W�����<���݆iΛ����p��t$k�E�5���_#�;e�m�h>��G��Ys?^�8=�����kƳ���/}
�5_�߲���Y��J���|}1eq��!M��B�ֿ\)�h�Z �E���JE�g���P*�(�p�N��!�1S#/��L���⚻�����M�^f�9v��#ܨ�9����t Χ��/��(Zd�bkذW:Q�u�}���#��
��}֢qc�3*��̩	���Af����di�}��������_���=��q�܉��b������B����L4�����F�\d��'�읪�%)�M돥���BG\.�4��z��uN|����:uπ��I��V�iO�Gu�Q�����'�m�u_y���C��ʒ� �}��;��~��R�#�j�����M�v��*����o ;i7��%:�7�Z��ɢq�/�w��-�s��o=� ��~���3x!�}�S��AO4�R���9��k^e���Y��e�?���+�m�}B��-�o���8�8����$Oīy��d�$V�s��y_��P������2��ǾQ<e����_��R�86�?,�����IK��jn
$���W��X��e�r3�.���9��:Is���y�x: wϟ
��?V�O��(������/G7�N�;s�]�e����خ��rr�G��=����k'd�ցU����95 A52�9��!�U�=�p�7�������v�ѻ��B�RE0߉E��������)}�G��gC|��[��s����7�_�����0uO����(��UeN���L�ĘM�/pU��~��TɤĄZr�Y1XTˑ����2�o���� Б��م�z��z�.ﱵ.�Ѳ�8V�Rz���g]	���
n�̟�;�qDŷ

����E,�r{0�d��E�#��d��(��R13��%��>��7�t�,��\�{R�n
*׬H��e^'�2ݱ�_�Γ��j�J����n�K�L�ͳg��mզ�����b0;|�#j�0�!ZoH�Fx[�5�˥����P��g�ɍ�!��]�K!D�%v����F4�nJu���)uӫ�<�q N�o�E|�I[�8 ��c��V�5���"c�t����Y�ȥ�8��F|�����͂�@m�$�e�����p�T���I�1�/�q�0����ᣬ��)�K$�4�!��g�Ӽr*����d�q��)ݔ�aa�9-E����4W�<��E�z����1*��6+��5b��K3%u��XPR(Z�p��H�E��`wI�4�u#o@($�=���٢�:=�N�{����p �H������~R�o	�\�! �?�%���,��d��2�d�nb�vű�Rް�hf�hi�Tu�y�"u�l�?j�̗���_B�=��е��{x9Ǩ�g���0�F!�b �2�A�~R [n��&'��ef������0١��knݤIUgySw*�j;��^�_x
��)����E�o��C�BooU.��n��<gN��{S���r�w�H��(I+%���}N�E]�\�&
}�%�G���p�9�h�Y}�G��~	�`3�d�A�IK'$���7�0a6�O-��VJ?�XB~�<�4%���Q�(�UO���|�l�੦Gu��a���%�A�����F@��AQ�pϕ�8c�陥MF2a�D�/��o>0Y�'�	��.�q%��sU�n��ݼ�uHѬ�=$̃$>��Vf���r����b#����jڗ�)ޮ��Ŗ¬�!I����?M#��>k�L�#BK+z�5k��N���&�i��W�
ŗ~��E0�24��/!钞��f��GثCkfc&����T��$�����V�YbQĚ8�wЖ�c<�P;���\l�8̚D�� �gZ]��M��(
~��._b�^J'� G�:j�COEX����;a��K����3,a�Aq��-�C�C�8���V�g��l��]�T��W劭�m��x����kP�2�+�<!�������q�I��?���"��+��-��wgs���o՛n�m��y��6D�<Z�)�,����3W���8�Wp���J�@�s�p��@��_�f��`��/�q	h�w��&-��]�^���/��(��Î��	��^�P�2R	ciC����|�{>/��j��Z�$�$��^=N��9�1��_T�=�����)�-VQ�x�eXL���M%%��ƿ��T䒇��=���w��b��fÇ;3�d5��C>�ds�0ېB��Ҁn��j59��K�]�N����0=����5���s'��`��'ٿ�0L�H~�<Q�!�^~9�l;Q�3��=1��_MO�2�<��i��H�bJ�ځ>j��m ��������7���'��>0T	+�2�X���1]:��x���ލ�Q	�?D@dPʚ_���|�1G}����p�	����B�Kx.oXv�<���<[�Z[٠>]m�e!����!�z�h�Po1���2좍ԻlE;����(.�L��[K:=S���Mo��WY:k�].2)8�<*�{� l2�ɮ$�y*2������~�%���ut`�[��������^����\�^xV R��2�A�P��D����ͱ��)U,'����0��Ko �j�WI��Y- �Xa�ʃ�5�Bg�2r�P����;L+��L<Ng��ʐa�]�%�_�2Mty��c%���Npݎu�����f�O%�R�wp3���1�!}����ȤZ�����>�������yW��]���K�E[��i�O��x7�z4���mmZT1�x,hQK�9����l�P��1�i��+j׀��'
���jH��a�1H� z
�Ne#��J��P���K���)��P�"\��PJ��|����H����Yb��]��nIqwDռ��V _���6(���C�,��b��d�Ao�E�!��j`d��-s6�B{(nP�e��A�U�|���c�S
!�|�vc�*RBZw
T~��V>(������3&:�PzK�zϕk��}w�`�W��8u�f&3s��� d��9��>�w�.��9˵�$Ϧ~�JV�JV�^^���g��)��cE��N;�Ab�I�_bf��E�kp ��;�b�p3�	t�I�X���&���*�7&>���!���^ȕ�e%�Ú<�����P�;�����F������đy7��TC�"W�h5��M*x��b�+sl��n�p:4>$[�żF��|,$ycb�zvQ���m��$���!�,m�sR��r��n?��E��+}'C2b��[<�$��^Ê7
�h:�(�&�F9�q�2V�R~��BeB��&�61Ar����js%Kp�6�G��H�d�Z��p^��0K%��������(�����arhzJ��B�a��=��%u;���( 9Ƙۮ�K���a�*���$I���-��j�ؗ��V�d*;��Y��cgl�O��ȩT���Fj�g®0Ԙ����z%��b���]����H'""X�����⃚|�g���&�]��n�����ta�����5�@�%K�k7�~44=x9[�Z���3C*!�T�h�U2���i8j��9�f�D�ۦ�n�%�,u�� \� �ffn���Lp��O��{|���5bp8�R(��@�?�u�7<�����^=˿��la0���V�ݏ)N��
�������yx���O3����4���4�T���&:�m���c�:�I��Dz����g3|�ꑬ}aA�e���'-'��M��X�͹7	.<�*��,"O����%�YZLo$�+�G1"*M���C��0��Eu�R!7�n�����;�YY�f2�J��>���sM��Cb8�i��s6��ᦐ�V�+�f��m�U^MK&�jP��g���1u!��6?s���[�ؒ����J�E�����1���_r��ݍG+�J2��"�E���Ը����O��Wqc� �\�-˺b�JV�����s�7�p+�V����1�ǪYM��*���S\��?�P�J%���~(�$�V�=B׼�8Dbh�ٰ<�^�/���$_(ss]]%�ZRG67��J�@�N��XŬ�жƪUu������翀l�z6����Öl����Vx�̬G
�K�R�nY,x���u#�Y��p�����"IC��Oj���o�;���I��{H�����G�D�;�9<׽z2�}���N�~�`��և������0x�}��Z�,E�E��F�9�Ջ�[���C����<G��A�{PM�� �gPw��ow6����q^+���GM�$���M�$2�E3��5������OKQ)�#�/y��N^ƚ����7ô����t��>�@^!ev�7���猸��ވ��*蕭����7�x�4�5D{���GK�.�6��q��}5`�s���_��ƙ)�c��+b�����Bĸ)�D,*dl6����.�W9�%9$��f���eh��oc$�{�����B�\9u�V�g��:��
wɴ[�u?���yћ (��^�K"8�Bzݍ����-i��'1��^gLѻs����o���4�0p�z��0{]Bi�F���D��ǳ�TɟW����MLoA�.�6�rz��F���|V�io���x#�� WxcS
7;���<?�̐\s��fw�Y�~V�[ђ����-=N���yBܛ��
��`�������W��^f���yX�tÍ�f}!\Į8_|$-�M�}es!W��{���ܸ��2P`ځDw�ʺp��$-=�h&!��,�-N�Xp�h���ɳ��帧@�+�]}���*H)�����ԋ7Y�N�9���BP�ݖǋoa��襬)0x��2�T��|��Γ7���3���9��sx�_M8���S}�$y��(��h���'z�c�Ԟ�&��_6�ݎ��o��g�ʁZڛ$T6��ѹ�,[�i��pƩO�f�Ţo�E
�X{��s�������[?>`Y� .d����/��[q��,�z�Q��'����cٴC��wN�y����K��эr�gF��F=�3��cx���'�s'h@;q�
�-X��6��1R�D~6ieD�4�5ؒ�6���z�x��?m:��ƛ M��2��af�:�z�xC����c�%��`V3��O��l�6�߯�|� �9��hDe#��6%B*2I��[��:Z������-�P���A_�V�3��������$��my�u�:A�y�gܶ�Ap��:V�#�&��)m;�k#�7f���Oɑt!���ȶ#6_���*+zA.2���z�ja<����nh#�]@84f�(\������#�k��_�y�I��np1����I��B�6����+m�0��UŰ�j���$�y���#��9�$�N^�8���B`=C�A-V�iy>g׈���GXmm8��ٌ2��GS�LM�4z[_>Ů��/��z:-����:� �:9����z��_4�����}˞�)���!6�Al��9./�9�$�Cǒ��a���_�M�a�"2t�.�w�Z<HJ��k����Y�Cj�%��������D���A\z@��En���+�����n������E���;&γ�5�.đ�vt��T���w,�K��6�<z��J�6��B��}�o)A�U����{��HI�D~�ۘ䐶��B�Ϲ���3Э�^�N��<2T��Qe!,�3�4�+��s���B�Dow(�L�p��»���*>Ю>i��7��e�Z����~��v���1�I�T*��e����T�_�=Î����|�����⊔3���2ζ���=��G�c��!ݻ.*����>A��z$���0c�8EɜK�K�:����Y���'��T�`��Qr�?�8�PIE��lt)�&��#�i�.��m�4ۅ�87V�NX���.�sZ4�� �ǰ�����oqCenw�7>�O�[�-��b�R�|�9�{�?kH�zl�']J�2��� X=�!�=v/@��:=� �<��JF��`|��+AK��+�c�.�V̚��7�e-b�y��a2gT$�R�1G��x�\7��Z`'�G�w��E7��ȳ��^P�Ԍ+���̎�9D1�-_�����Bgw�\'�&�5�(�~��g��P�rXd'0#�L�ϼ��Sc�(�q��2Csȷ&5���`%O$����I7�D6��\��5b�k�Yq�<Ѩ�t��qjޤOk��U+�MXqf�������������������m����1/�_0�23�n��Hs���L�[�#?P1�T&n�3�����kL�qe��0E��G�D|����!y6�ீa��`^,��jö��Jt!�ǈ���VQ�3��x�(�_dd��:�9K��k�6�EO}��t]�&p1���MX�V0c��J'C�bLpkɮ���]hQ>t>�d�}ݸ�jS4��k	��A����Ʉ^g�����a��Q��d�}���S��'�$��LO%�>#9�|����L�ٹ%�<.`��2�a_��w��1ޙp��g��X��aq,U\ M�����SD$Y�>��Դ@	�*&���>#RO3��|u��9�E1�nYt���@�q&�hk/
=Pt3ؾ�ue�9��,c���:<�.��iB�6�f,�<�6����y�Ī�S���K��_����X�#f.ƨI��l����Tg`�5�0?z����Z6N�{fuB���L�ӳ��UGn��e��y��Ad�!:�M|�)R��Q��P�o��nH��?�^$�/��۴7P��'��w�*�px�}!1a"�-O��ntD�ˣĀq���^^��<��9�VD$hF���JzQ�Io��g�ۂ�%	��B|1{��S{�c��(`�&�$Qnu�k�AO>R1�v��c|�T�k���7�~\&�l�q摺�����E)�@�����`���,Iqz�N�w����%-b� �e��](�<M��/��H�_K�]���!���@�V���W� X�+����χ*��w�'@zJ�R5s���.A�v�L�e�i��o[��8�7[h��M1�|�;���[`<�N^��٭��>ݑCy�#��6""7�ڛ���-/7U��L9˯� Pl��~%�6�FD���zA� 5p�:{����l�
��Tf*;�m����eS��z�'�CI�#Hd���@��K�x���\)q���\x:��l�TP�����XJV�z�K���ȵ��K��]s�zt9E�r�D�P���G�;W��>��2�i[b��1S)r��x���)�C��Տ?�������K���Ct<��³�a�������TV�	���z�.۝.u�o���R$)��[k��"Tb�+N"���	nE���N� Y�Y����nJwF�P��B)�/\a��T��������\�,5�>��B9�5(I��<�	��ˇ�Xi�|�'�����G8��~�o����o�S1Б�E�h��+�5�O��d�)��"��U���3�_K������c[ϸ�gd*@J޼�eY�jV%`������?)t��,���O@���-�R��-���N��3у��Z60���"|�z��я�Jc�P��_�+/�zRڱ�XA��{Y��{z�n���6z��D��'���jx��>�"�\�0�sG�Q�a�Ϙ�/p��S5�}�����S�\��g�=O�cD<�i��k���p�pE�1����RK�p+*�pײ�E�;U�+:�^�o�h�SFcE�>�h����*�Z��wP2l�	���UʳU]P����@w�t����P8�k��ߊ����s U�^g���Vc"��n7��S�_v@���li+SV���h�W��y���17��U�ر��0Dz�K�zeyF/6j�!��ڲ�d��+T1����!����_r��o��`�����%)����m%j��N�6K�J���v��+/v���G��YDl�F��&P���N=�E���=�@g���%%O��q�;����*�O�?ƍW"��.I���X�{#��w/�r��å,c6Gi'xA�UԢHL�0�`!w����:84=à[i�b�8M�ˡ�zh��l���G�48�#$3�� ��/��Gȗ�������nʈ����̔eE�{dTW��]Zմ�Q��-�!�(C�(`�힨u$�<�2=�s��N�O3{e�Nޫ�C��TwV-��6xR����Y9b)���j�&q��A�V�&�:��`�ý���m?8
u��B!���)t�m�I$�6G����j��c"Gh��������t2�>�������aƥ���nQGK��e%.G���rR?���i���R��MoP��X��p���]	z��pUŰz�5Wҫ�:箶�����
�/�=M �W���}�!o�s��^8}�KeGp��jz|m��*qtf�,���*�Y�8I̟R������`
E��C��RT��$SS�D���IP�0/��V�L����'���Sc�~�η��*�����g	����l��{w�T��v��YA?��Up��P+җc� n����ח�u�U�D��H=>���۲S��5���Å�N�a
��`b�g-��}=^�4��x��H��a֗f�b�\�쉤����w�E��� {3׉�=!�d$�>�{P>��`�4�dG1c?^���/篹 ��|r��/��Up�B*��ڍz@mȚ�ť����d�Zi���F��`�E)Uק�Q�d�(�C�ѫ_�6#�@���f����χ�nٞ����@%�	���Sd
b5SDa����J����;*�D��y�#B�2:̟!�������k�8��e:n�)�8��>�B �=�r�E<aF_3�c�=�j�u�5������!ڐ:��S���q�*w0�|A(&9@{�=��r�vߨ�rE7��/�-�5�$E�R�=,���� ��Mm�ܷ#����+կ�[�+�D��,^+�5S�2tc�#f�PV%���=�|�I��e7PRn���|����5llj-0��ׅ,XC��սp-��L4	�El�U^c��R����H�P^~�H��@S ����;�����6�7ܭ`�^��PRJ�:5�h]��x��	3-�4G̻���ݿ�֕��/���?ْ�
�"��s�L���%+z��:�#b1c֢���F�#��1-at����]�%�w:@Ґ���L呬)�1��B�!�8�|@�~i�_���?E�9�N��͢��&brgʩU�^y�ã���j��0�16� �:\ �	¶��:��Q`��E�ݞg���9�Iv�JO!��=��И���Dml�kΆ���G��@b=?�=i#�?^G�w+�M���m�eR��*
��<)�{��{`*>^)�u�蠷zZ,�bG�������+qzT;S�y�s3�uq4�ES-"D�kr�`��0.%�K�c>�����*�H��ݳ��j��q��tˋF���H�Ei,�����M�1g��[�D�������BU�|3�(^�U���!�d���d�8�:'S"q|Uޘ��?�|U�oL�� �m�����[�A���*���Z���[A:u	�L��	�F��C���~�A��||��ȭo+�>{.�����i2�˻A�N�`r���JH'`����I3>;��%U�[�e@�6ӥ�?;��Ox��%k��#�*���goc��a�����j�_��4� ��~�������� �o������xѻ�k�Ğ6���|}�t}{��D��O���jp?Q������@�T�6�=ت�ay�z�;�b y˳嶧�o�M�Im�ȃ�s�G����h�{t).�Pv�f��?�"��@�d]��L�����?��곰��a�y.E,�\ �r��_��/������I?k��Äo��U����p������$k��
�����[f�?���VL�(�`�hHzH�J�]��������7�f�d�O����h���
1�Nl_�����Ȥ{�]k������)���鰃���E�b�͑�w����כ�d:�Z�:� XfY>��JC��v�0�1zގ�_wv Sm��i�^E]�~T��vul%� �`Հ^����[mCi���P��h{9��HC����zvV����G+M�ꃁdHa�t��t@a\G�(�!"�hT|����j�ITH,q��ߜaF� v$oa�57W�`�Z���E�5y��I���79������"��A0�΀k�s�f �Me��.s�v�Ƹ&�Rj(�̋hKI�t�H�A���r��z�Iu��JZ��P*���x4�U�
��h[Ǟ�*��ĵ��.T.LUaEÆ��K'����w�e��-�/����6v����WxH����-9��{�ZV͡�����r�T�����{�JD�9���1�a�!�2�ͣ��	&��V�X�jK�ӟ;X�:v�M�z�?)�%,�{�ɻ9�ü�����e�>ӻ�Ө�x�?���X��8��0Q�Bս'1��&�z�7�G6Q��֫�r&�1u�O/��wy[���M�i��}�s4KVW�a��e��1j�*7���yQu�%��d�Oң�}���n�p��� �8��� �H���&&���8D�&:n`k���%7ڃ��?4��/
�C*AE��J�V�]��ƈ����(=���H���"���ެ� 6�rk�9����-}���ۉ��܏�&�W�<�T1M�޽\�8vmc�:]��7'�ƪ�g��y��7'5�z���Qin�.=�讂����$�K�K)u�]b�++1R$9}2H���ܕ�j���&����?*��m����8��,>n��fSG�~n%�4)�	~,}�Z��0��8UE�	��ksg�.=�!
u@�5�����ޟ޴�O)���W�f��@2�t�MK�_�j�c�N��4�A������};`���P� f���u���R��H2T��I��΃'19�����M����nsc?0v�F[��jc�q _-�ڂ���W��zeY��K����"�N4V�]����J�D��(9�&���`��Q@��FG qy��[£V�R�-�Տ�v�����ޝm�1���AX�_��%���22	�w��
W�(\4��꭭����0�m@����aV3߇<� �:���k���*����o�5���|:�+��&��[�4UWP:+G�U��+`��%iN�W?���K��!I�� �����,�G^s���+:�=vrW`Xna����DD��r�+�����}V���jg�`z�a�s�_%%TSe���	�m�<z*<��E�HAY�FF��	wC �d���!g�,��m,f���HwtR׵�m��r����?��'h�V�WtSŤו�̤T���F�ܥ���'��1-���Ǽ������N�]���S�۩Gkq�j
��(��������`۴i*�X0����W�a_�o }�:"j��ꪽ�޷4ʧ�Kj~ �^�:﬊�[���*�Ce�E�o1gW��K����h��R������+|=3��3����]:�Hc�G5��J�.�ܘ�Pp�tӨNo|-|�B1}�+�-��$�rPr���%M��-Vឧ��o�PIv�ps��G���@"Sv�K�&�/rNµf�M&4i��¯��V��V�%kL�y(�>�t���Y������:�#_�]󌣷N7f�ٚ �]v��b��h�%�-e�^)+B�6�
EB�to����C�:�v��z����^Z�ܧ�H!I��/�>!�=��f��u�]������,�a�(U��ؼ雤������,&�גBpM�4���B���Zc�lG�2`��8��SnF�m�쩹1�WR�rғ�e���-!A�h��K��N0�jF����n�`ߪfd`�G���d��v3����Z)�/p%#�� �/��+��o���'Iz�)y�0b�#f傈��ka�J:923��r�%��Xo\�$IբPq���erߑ��������`bP�e8��r�i��ܖ��>������	����9V�
�pY{����{rn����Pts�0IX�m��=z/�I�2H��{�V�V�]ⱁE��'+곖-8�A<�h�J<�$��-��Ik{OS�_����fItpF�cm��&^"����JP��(�8Z��K<�[�)ů�ǝ���Ys(]�|���]R]��҇W�ާ��Х�`!���I��c�s���F׺�ٓ�)���m�d0�ǌ|�+��/����j�n܊��z=�1f���­G�hA���~I/l�rh���^|��%5�ԯ�֔��I~r�/KqEw��.�e���|d�.�L���Tg1�H���7�e��F.�9�����:�/�7�('���@"�� 8���8#�]O%�܈�M�����3�^�+�2� �i,�����A�� &��6kC�/r+���'�5?1V�媔�������P�~0.�����|��X7 ����8�� Wڮ��w	�={V8���۾x�m�����gY����_�i>�1���5dZ�{�74=dD[�]�ss�vc�i������o�4���RM��,�c��!�"`��8�GIbe_'��A�܏��.D.v����3@��Gc4{����m��*rZ&� �
�jP��}#��r��3��({<��c��i��8wr���ʶ����.�RN�s�)�x�\~G��W<�9TX#.�EU�W�|v��d�(��9z��RuLg��&6��������ŌK�T�V·>����Փ��P/��/��<+`��M��E�vo����i:C5du8���/��+���X��ڿ�+(�!̗{2]6�m󓴼���k;.�7��+��G��q���e��oM���4�k�n�u<It�X�peB[[g3��JG���燲A��n�Q��������\Ey���2|0�%���,L��X���'�wn��'�G�y�:�ss��S�o��b/;Ly�	6�χ,������rm�Ɯi�_��|ٍ�ς������w��Ʃl�ڊ� �C��x�NI�6�i��ʃa, ��;���ޘ�VQ�e~ϼ}�AU�ӄ�k���r?W@ {�!���b �bAb 7��֕�&���[��&g�$ J7�����_+�DRn(�a�(�T@Yz(�����>��9+K����\Y���	���dS�M��P�h#o��!֋YF*�p'^���5��ț�&�}g��]�Pc�[�i��:^E2�O���FX��N�cM�@��Tr��0�����IX��Lb���qG6�� �ɪz�r;ڐ�!�m
�ե�&�Wy<�F*�����6�!"�C��R攣�`D��h��`)���yQ"c��Љ�l�"��]�F�Jz���C��+�.�/�6r�L�z:��=6��˞���>��\1&���Nh�5��>wY�_��\'��t\[��1���a�}Z^*�m����6�v��} r�v;�ކ�^�U��F���/\�̿���
�a%��OlY:��j� ׉m�q�#���^����8
�-�AZI�1\ݟ�UL�<�s|5e��<�[$����r���"���r#��PY�� P"��f��V}=�)���) �KV__ްO����])S��h��L88�����j�h3Շ�*�������]�|�uԨ��![^��	)�	�ܨƃ�g�1R��M�:)��7+�E�4[b�#x�|`j��D�S�j��}��Ϳd�p6Y)��q�2�C�JX�7���:.dkdA,]דf����x�s�˰p&MPfSǐ�����.suy�4)9Y�c2m��I�����1g��J:^5'�n�!Ai��b�9�`�%!O#��Eyg���M�`�.ħ���\qen�(fo�Ϯ<���&iR[u-�R��\��F�!�a�݄mm��d<���D�罴w�&^+^j
���iK-=�#R����υ,��ȶ���\����C-������+\M����V��El�jH��S�79؋9%���:�buڐ����BU,X~=.�#��re/��H�5U���|�:�ۡ�I�c��|�A#0�Bo� W���8c"M��M����@�FGٲ��}�@�qj��J&����O�PY�n����#0���k�Y�LE���8e'� ��3�-���UiN��]1�2�\�(��̊lF���@1�>N��W
��#QB�\x3nR��W���Rʗ~��i��C���-mS�FDa��ڡ�n	f���k:��I�~�wq�ޖw���񾍈1Ƅ,,q'��5é�6�mNM�H&2@�f�#BOӊ̐̃�*{_��GΌA���.�m���\�l&��f��WA��z-c�6s��Wc�D�Zs���M�C�XG�S���e�dqC`��t�0yfD�ZǴrܴ{8@i��?ݣ����Ԭܚ��}���;C ��1�O��b�պ�W��O�uܫ:�{�+<&�v��\���~c(�#��Ki}����K��êT0յUk�ޥ���ݢ�:�#����̚�Cb�� ,/�
h"����oV#\���\��Ъ�ɍ��e�@��K�Q�>���-yCd��,)�[��-�ŐN2�uR�y!zC4h�e�)vH&/ENL�Q�b�����$%�U�u�D}��J�O��% M����6)���W^Mp/k�Fl��#���p�n� ��p��t�����d)} ��G�{�s%,-�J<�`E��a��ܳ=(�k�@N���C�{/�S��B���H���"�&��sʣ�a����HX���bwc�����Jf>�?h9��dz�p] 7��ЅqBD�It��{&��$h��~c��T���"<\���6U�ק���7~� ��������� o���a7r��r:��'4�y�W���&j������C[�\��Y��_Uh�J�T��H-�L�� j�c5'� ��D�P����$������S�I���;�\D����!-p���=$��Ne�\�j����u��״���I�ã��û{}�M^''$+�*���FU/�	�!�)!�q���4�p���U���}�ڂjP�|�]/�p \��ݙ�3!<����oV�ΐ)z}9o�H,@)p�5pZ�F�v�-`B>Z��1�Ԍ�>�cįw� I9֐%\�3�%�6�Q����R* ��إnt�����02_��vT#�b�%&K��Cz�a���1�kG]�|�1��f�X���9z��dq���V����C��I .pO�gDV�i�����/S�����'07<�.��+�Kl(u[&Wh�@Y%����-�GrRt��kx�WU�����۫�.��c?��s����k�xZ��[��5+��m�K{�K(8f��͡uU����65,��K�h���)Ѣ{J��Crb8(����s�Z~�ÿ�bCo0" ݹg�	k�̼���xh
����EL:�W>7��������Hiz�Ab��"���.DiȐ���j�Ȕ��� �[����,I�E��#xh"j�	[�3��4�=ƀ���9�$�/C����n�8��4�/Z�tq���hݶy�a�S('���FT;�z��KK	 �s��9N�3"�Q+m$���],�2��8 V�*� ����S阄5kd�O�$㸍�([��	�낸o8��R/���=���Z��FI��H������f-�t>2���a�C~��L��
� q�:�l,l��V-�IKٿNI��dQ��ׇs%��9�T�Y�d���*�2ѻ�����3�+[��l��1��!�d1$7���mثL2f�0��Ń�[�٧L����e��3��<I��{��N��E�k/������7�(3ХXӁ0�S��y���Y1;���@���e5~��I�=�<Ή�N�#��d�j���O����M����R܇��,�]k�@FO �?'+ j&�k��Ҽ)%�#r6P���n������������i�@=]Չy����;�������b@uzL�
��F�����f�X����%����VU�GuEҚy�12M'rU���ʽ9$.�Z� �֍���0nf��]�,�=� ���0�Es���_�z��7~�����.nk����Wd/9�� ��y�e����dh�1��-�n� ���W��\Т̣K�Dt���~���h/CZy�AM¿#��u��eV��Lqqi9@����6�O���Ɩ^vK��D�d���>BdDRx�����-��3xq�̑B;���@���"�{�cUhqLN���8*��	N�m	�RS(K����h͇�S���m����iUU�TZ��
��D�[)2��oh���^0�~wH�D ̾��6+|�+��1{M�����xA��hB\W�/ۄ$���q��.�����,�'̩-����*����M�uuwMn�B���(e�aܯ�[�5ܟmw�6_�e(��χ�1���6'>Y���Z�W�G�F+��ٹtF������<(�Y[+���'�o�Z*��gk�fȨ���t�!���̀� HE�[�����D~�Q ˂+ӻ��	�{��GLΟ��_%2�ΓP�K��?%ӝ�����#{|�/�%����T�e���\�� t��S�t��ƌ"4�	I憅�ԤȊ��Y*D�4��(���� Gm�F�� 1u�]��4��E�6��@C��L߲�,Eb�Pۣ�ϖ
Yǭ���ͽ�!)�*�0��uV�D?V�6���l5*�C�BV��G��kDx���a�|)����O3�"ׂ�����琭t6�bG[��
.�E����+w�k����|�7np��Z�*^��g���D1#	�&��]p�WK�, ��~w�?b�N]��C��	��@z�6��A�����m%g��l7����y��b��ܩ�	>쓛����Rr���c�zY ٖ}��¨�
C�'�%䣰��g3m�L�U�![�KnƜqt�ۂ3C���%j�ʋx��;��o��e��wxk�9�����-I��wP���X�F��ӈ�1�RXZ.z^�Y�CU;�NnG:��^�c�Ѭ�Ң�%,����)����l�,�Fg\/���]-�3��ԫ\aeN�>�]1��JK�t�XV>�E���z�L2�@�B�6LĹ�;4��aW������R,�
�6��:K��~����@�����z�U:�<<kϸ�t;_i��Qi�0�v ���d��9l�k'�%.�	�MI��Ѫ����6��"�Y�����2�S?d�0w�.��EϯX"E��z��X��"�H�������_����A�!�!j-vV{a�~*s7p1>�3�ڻ��8��驅iW?�v]R�'1�s�߫/� {����D�KJ��0z�m;ǙmE/d��Z�6H�)��w�#2^/�<z���p�{��+��e1������,�I4"��%	�j'�@���$�4bt���ݩV���
�9��PyPd7s/t���.������-"����ǂ8�����c<͝��1v��Ƅ�^��s������4��Q_!��= �\�nX�NzlU��i.����C[wbN��첶�OC״^��80��gXY��7s��'���4����c���c�o�nJ�?��H�E0Mz~�)���;��?��F`b�|2�!�'1)e�D��c����7\@�g#���ҙ���S�A6u#��_zO��$��%B󯹇@�M�K��:1��=�-� +O���L��q�"iyI�oq5�:�j����e���̅�S�o���U:��O�~�X�lQ��b�կ��Dlo�����ʲBpN8R��j�"?|�Zb�]��ϻ#a@�d�NP�7* 
��ާ�O�=Ui����y�q�sh�Fm!��ɛ֙��>h�jQ6�SQ���[YlRy�lO`_\��d��S��J#w͗�DWF��Oȿ|*�$�iF)�.Z��	 N��n��b�r��/��@����[w�g��\9���@$���4�Y���F=X\��`u��5ES�݈h�N�A��07$����!pߞS�L��>��+-��������a2�:%��Ӻ~)�j' ��H }ru�"�$�ٮ�;�[)�{ׄ1_�혃�<b4r�'r�L��4�>�%���ǽ���f���Ӡ��%��E��!�AX=Y/ַ݈V�k�/�J"�}$��➄0���_��"}!`]?�8``��b�Zy����z=tx�`@�>� �.��W<�ov��yҋ���5���C���a�uΖ|�6��\�� �w�$����T�j�?Hx���Yc��F�`����؏�9��tP��$ȎU C@=r,��*v�A׀r�et�}ؽ6�o"��uo+%#�]ިQ�_�ɐ� Ȏ̉=Z��O˶�ڛk�I#�F<v-)�e����R��T���M��{��ʞk��t�b��+�֨H��ؔ"N9ھ|ּKR]��$���t]J�B�i������VЗ��f�f�M�=�x�4�$W,e�<gKNE�,x7�h�_|mlS�� �&*�5SÆ���;����P�s�䓦���A[�s_��y�;�����:�ͥFt�Y��י�~��[e��	F���%C�ΐ���G�B�)l(�x�����t���f䟸�`E��F��ĐW�8���gUXf��������&0��-^���6H�C� �ŭ]�b\��&J������:���M2����Z�zrrXiȺ΍h��^<.AI��X���2XÆHHU���4<���l�0BT��H("k�pW
Ѝؚ��nqV�`��鱯/��XY�jπG�XFv`�*^tFe�rzR��e�ѿUo�aP˟AZ�]�� �<v�����yC�GS*��RbV��N��\THh ��x��E	y��E�-��|��_�)Kg��W�
;��Y��U-�ㅜ*��k^���n�&��3�(|��8���x�����p�i-�{,����F}�\ ��J�L�����?ʔ Ĕ��&7��˖^q�1��-0�Y5�w !�R���H���[�V
Uʰ��U�,iI>�%����q���^L&HB'�Om�[mN�ڨ*���	��Y����v�z�Q*�z�L������Z�i��u�j��4;d�|����@�d�fɏ���ns�6��D�A@_ؼL�NؑyrU�������`{t��;+(aQ&��VW�d�NǼ�$��"-������h���CR3!��JY_AϮ�2�h�pc�g�J*&�%;M(��T˃�Q��|~�3�ďl]ߧ�'�7��\��U�f��/��j!�f�1yg���n�b�mF>Ʋ��2ӫ;s�Ro�%��pq<Q!N6S�n�b`�5��V�䬅%(7���Z7��y=��=�P<����ie�γJ�b�%TtI�?���,q�(	�n��T�XfWK���%�y���E�m�S��@�'�|��`ݠ�f��-�,����\�E�^���I)D���=���:5B�z�*;���}�ӥ+_J�u�rv���"y�4x	ja��V=�$HL-���t�0�PT�ny��-��ݱ�z��J�J��;ˬ�R��¼;5�̤�$ Bc zT��bVo�8�j�u���E�0��{*��<��/�n&P���
��ꗑ*qr�W��V�:��;=Ə������'@�K�(�cW�qL�1����]�k��m�3�FMkXuM6	�?ԁY-1S�Ht��P�F�+�I�tu��EI<P�[<��������_ ��.�n&SLaF�tW�=o8���ž��s��5O��~�R��������\�W��m�#}@N�ڨe�����f&��8�/���%��GB��SbA�B����D��g��s䦜bO^�ސº(���+��Y���Of�34S$<q�G�F��~�aؕ��Cu��$�GL�@����ᘐ���A��� ���0���Woe�7�R�xݵ��3=�%'�29�8�[S�� �v4)�s��o�L�i=���p�1Ǽ<�gzV�~��(W�B�Ԧe����na��,z|N�i�M�ScT�F�6����,�f��e�H���i��e>�$ă{�$h
�4�[{�A��#s��h&���e1\�yN��D� �b@#W��l���m����ed.������îZV_�3C-nu#""Q�h���k +!?U}$�x.G�����)~�v�,Q�p�g���s�U��cK׀�[+6vo����X�'K�D���i'�ZN�m{��>��¯Sgѱ:0,5T[�@$3$k���K��@:�0j����Z���
8i<*�t�\����Si�S�.�u���10��f�[w�Lm�יuv��dQ�������ZI����3���{�)P��S��.���՟��#���5�y�����f)������|BEl
�L�+X#���]-��R��V����}Å��`�[�>�B�ͦ�F�	�K;X;j1b4�I��d��tX FmV�<�j�x@�V��uRz=�>Ļ#щW<++_�D�r��F�E�T"*M��lX��&o�)�����E��*b��9��+R���-pwm��T��D����
���>�W	��yŬ�B����'Z�Β���#�x�m1ҭ��3����%̾3�G ��8mOmL+ï����:���p=�p�:Y����1�B|���|*�F��ǖ*��%��Z����e����ިx�|����~��[ʶ�/m|}�l��
Qb�$.�韰4OQ�D��Eْ ��n� �=�6��ך/<`n!9��h��ԝo��� ޒ+#v�J�[�y��/�@�أ<��>i����b�{��뮺���h �#�sJ����.��H�>_d/������� �^�z�=m��_��������-�k�(	��7�jݘdgŉ��{�+rw��O�]L�=[}��b6w�_��$�^��e���7��67�XCf��d�Vo��P�Ok��5��FЎ��n���I��4�u���ŭ,7�ۀ�bpY�;l~�׀)s�ݎ���g
�O�b��w��R=q<kAsض��ي���s4(��
�7��f�80���߼3��Ūa��ښ31����gҾ�G�C퐵�b�Vt�͓p���}��P16��@��W�6M#�_5�)^&�6^�kA�B��p��"C�
�e],�O�%����w�T�ׄ�m0dnv�"������p�ޢ����c��<?�Ä����8W[�T���V�9(z�&�!3_R/��	Ёψb��s\d�㰪��8��W��9h�V	��_(���N`�{�nTϮ�8�����P&�ЁJ5��`_k��$�~�ZL=�q�5v=�
����@A"�A�8N�Mr�J 9��e]ӆ��?�[8�$�n�{s����Pt�?K���T$���S0ThҮ�V'�N��訛yD��/��ӻ�[���&no«���c�cȅ���w�aý��o�����ѿ�Pa�R��c�����,����H̔5�_E�@Ȝ$��U�p�]&����e��B�L@Ĕs���s�Y�nB�8_c��.�hE��-8$�`\#w`�0Gт��΀�l�Ip��ր%mv�q�7����P��O��r�df�6��=�4 �hh�E�ӊ��d�u��K����r����e��*��p(J&�up�D��|�/vV��h�!6�?9�«��2�a�&�G_Ғ��_{;D���|�.��E�(_tŲ�k�/MB��g�`����~�h�"���[TP83�5��H���"0�ˈԽ̰/���L����ވ�H�oީJ�7:!�O�ܿ���FD.�ʊU����n�8ނ��;�7�{ST�|U��,��0<0@p��ɳM@�.Y��G��9��R�^���|V���ͳO6 ���ң˺C�5[^��;��j�6r�������\������ ��t�PA6Bak#�a������S6�X�x��5���?�`e$�t��N�G��Q�##euF�{�~�W��HVF���t�7���&׾�(��(��g��%1��q0ki��_��� +PE]v �FUi�Uz��O�Q�6�k����c��s�[���n�b��S�G��#`n���&~Fh]��d�I2B�љ�y�s�R�.Z�['e=�:N�����Ζ�Ă�}S��Jy8,P_���N:��.{�Dz�$
/l�lʎ/�����A����˲hOsh[�� �ˋj�B����sO�幂��}5V�o��>�a�
�)�ፉ6h��DX?��Te��k����B\T��M�F�H�hÐˣ}c5B}Q	�wLd�v�2�kӖ
S&-��#���q匢�ð|�ux?*�t�U<����"�5:'�9�^e�������Z��,+�Ήɭ��7�r�L�hL�F��9���[	����pI�6����:����D�ŰB�]��J�E���,}�Ə�"�nO���@06c�V��60���l�N�T��Үm;/�j�/�ϙ-�h�t���u��me]��>����W`��5[c�w]]�Cp1����g��o�B��_�9�?�5�$g�n7�ǘl�N�����j��9SE�t�P�Cf������U�[�'K7��Ԫŭhoc�0������X��Z�����I4��V$�
�������_ۭ��n��`v��i��>F�C�$;`6�KWA���k����B^���z��#�=H�5}�����K��L%YFd�6IW��+���r��+�����"���#!\�V*�"����W,������2���23�Z����L>*��[�\��� �E������R�������~^s��l�����A(����RB�T߲�g+������}0�n��z6�OPБ�Ս��p��f���oZe�B͇
�2�4�A�-�������7�����i��p���rF�p�g~�,�����l��Q`ׇ�����<D���q7"cz��QD��&�n�¤��
�����<�EFן�z%��z��}�����.�?�2�eB�:q�L��6��$����z��y���ͧU����$2
��8��� ~�OBZ�_���9����Y�̶�������6$&~&�F ��|��p[�( n�9>Ɖ�)�����l�޺J�&hkuB�?����h=�;#V2��~��d?���(�0��IAjj��k����:&}��l�1���w��\"Z��	';Z�W3b�#�\]AZ��b�_ټ�1�2�f��(��Ǿ�Og���'}v�n�)	C�/*B��$�ۙk��ȣ��E�� �O�E�ل=�~���~9>��5K�m��~�B�(n"p�+�QA��=�bB�,��H�wN�9���耇�� �r9L�\:�����ڞ��P�P�Ѓc�3���n{ȧ<��Wp蟅;�7�)ϧ"��`�?��t}ٰ�%���9�l� �s���Z[유�W}�^X�D)ᙝk�U���FRm��+i����)����D!�R(��n�F�7�L��+u��5�7pP~6��e��(͑��O�����WP�X�p�pھ�w�u��*������Q�0:�sb3���^7eU\�Zӓ!��;?�1=ca�2����hjnc��xj��'�>R� :�����.��.?�xz1[,���7'����������0n�M����<6~�����Qu�v.%���sl�[LH�K����1^8��'��3�;��-�"u�����:i�w�(��m�-�h��^�-ž2&A+��׎6����*|� ��� �}�x;O�\���37�M�	��[�V)��jĎjߩX��v�)@XG�tdYu�|�C�'X����9�;��<y���jU;X~�诊o�Y\'hE�ic#͉	��Jo��XHy��ت���ݏ�~1�ɉc��(��<��r��V�B�MoK�?����؈����뎷��p��x4l��g������>��}��rP�#��)�4������Fr�f91A��Cx���<��H����R��;93��B��0�j9gFP�)?�ݸ�������B���*[��o�"�	u�>�K��f*�k�e��{I���]�n�f" ����F���n}�+^��-Օ	����->��S��Y���US��i�����(�]��,�u���΅A�Cy+����������%�&�i�Qw�c,�D��S3a�n���v�ai�`X��Gģ/�E�s�~q�@��bn)VGBf�}֜���ȡ\�B��X�%�ܭVvA�Y��/�Xӈ���9�;/��)�� ��[�cT���R��`�iKxdN�c���c�WV��{9Kh>	H��9��3�tQ���M6�@�����djӃx#�߻��$o�,��{:��Q����~h\`/�s,�p:��(^gr=���k�G�

5���Yplh���R�'v��M�!~H�"�Eb��	�#�\��`��J���}OφG�g~Srp�Ơ��bM~R�/�6��<Д�b>�E5�&��^��o��'���3�_��l\��I�|�'���}�m7Z���D����tJ�760��r��M�Xbvh��q��f�"b�tTk�4e��$��J#N��@�HHz$��{�#0V�.�HI�.����C�����S�q�X��VmE�5M����ٚ���+�S��(����ס�%0�z���(@^������K�
��	k��|�T�#$��#_ͨ~[�c��Jj:A�^"���8X/1��q߽�m�T�j�w��09�=o5�~���^���_��ə��+��ꗀ#a/�-����p�o��dq�m�����?B	K�ov��~=�+<a��$�����s~Խ�`�X�����rC]�U�zhH�5��=��ʶ��m���f�	5$��o�-+�z��W�dk}u%�:eN��������i���_3`[�.��[�U���x��[y��؆�)�+B�r3��b"�1
�Ez�L���I�:�Lڒ��$�$YJt,2��#�	fę��Q1v@O�|������L.g��!����?��t�����.�)a����X�Lخ"W�$��������[�ח�¥ؗ��e*́6�xV7���i���,D[����-V�D���γ[�ɿ1��4�1��Ģ�`�&���;����V�A^��X�ȟ)� ��~�_�x��	z� ~�Z�95�3�P]���ʖAF	D��XC�I�I�-5�G�����̬�]�n1[��U�Pk���"n��Oi���m��r������x� ����("n �/h�Ku0.JS8;z]�z%k�j(@�^�
�&�������5pB�����~�C���.B��wDO���
��½mD"7�m�c�� �y�x8�lh�̕�4 q���?�3}�Bj��T��ICjs@X�����N@Yq3v���n]L��,�40x=}���������˿߼��a^2u��6��jxE#E��1N�pg�*d�n��~�pd���o6>��ef��{Ը���\�P'�kS��RE���B־�� `'���������Pd��|�Vp�}-~�C������(!�pP�G�QL^0�4¬�m&/�[Vb�B�!�٢����ډ�0M�F��F�Dm~��APS���E9���%+\7����`�>AG��Z��f�E� ]�aHQI� 0���E��s�W�r�M�8=_�5��6ҩ��9��p��$��?�
T��7�h��˚%b������+�π~_��t��"�+�A�=��8�*�M�W<j�GxW}��D[������EN���y:�W�(�A�h���:��(�(����1t65\��鑞����m*x��~�-���t��4��3�&L�n5�{���D�'�Tg�&��ZF�`i�)���NF@�N��Y��c���"�w�]@~�߲#M+~�~.>#V��;�z�?
hF#���5�4EM�&u��}#M�����ŕ����7^���`Wq8���rz�Q8���P�3p��&63,�SE=) eq��X��tM��.-#܊��\��������-�%J) }����͍YM���e�8���mUO�6�/��t����n��5�%ˡahec�C�K��,�4�֠ߝ�x�y��d
��-�L��R2ʁ=����8߲������kI��/�A*Y^��KbY��%�"�4�W!sb>W�k��s�_zr=D��c�:�'z�O�7H`�#�Dj����>�	��K��O7
7�P+�h�{�����n��"�H�t�G�֊�6W�RA�v�I��,��&�*[r-2�FrOH����kB\Κ��(K0����7Z1Xh|�f���� C��`&�jZ)zMV(=n\��"8�Ƭ'�ɽ(G��9��t�����3nn��^�+Hد�T)	��Ȱ1����9�#�B�����T�(c�H�5���k8����/g� -�1F�o^)�DQ�aR�VO�0$��Ř�rI��h
93~���m1t��OԄ�=���-�2�=2y�u*�b��d��mv>�:�����17�� �X�%��QH���p�ڌ=暽v`�$�TVTI�����XӤ9a����c�̕�#%�:8���/6(B���X|��s��i1�w�8�0�����6�6<Y
�j�iLǅ�����i�̆�4��A�e��:�Z.��9Tr(?���A:*��1�o�
k+jz���U�]��X4��֟h��QJS���:Dw3;��������y��G�C��E?-U���G#H\���i��&`�)����0δf�1��rb��o���nn@��D\9O,w��'��>����`��)��1Y����<p����'��yMb���i�,��w�N�^]E`��?֊m� �.d%y!�+��1�J�(�i�����r��n�.�+�fBSdk�^&��U=�vŝ��D��x�N�\����G�f!�"M�@nr�U�ǎX��"�=H���@�_�<�'����cc��|�}�dd/]�ͦ}�F�X���(����8*��� �L�H{`f\k��xh�=� $W�hK~פ��m�Roi����4��X�˯��6�R�Vu�C�k)�%q�a�,`���9ȼ%+���Yf�AB��#�Y�O7�/���a���H����=hA�����58�$���79�@}fG��=d f�X���,O5P'��H�M���dK`�$�q����C5� �5S�:]s�x1i[�u���r���^N.d���z=XN7U��E�!���֟M�O ���B��ؔ��:h/u��r�hAe�c
zC�
"@����)�Hi�M���2�:>_�FO/�#�1	Q����N�W ��֙��;=�����`�w7W}��|V�uB��7	��9�+�V��G>#@&�׳�+~ga���a��׬V%]?�}��h��
���RU%u�l>�TN�A׼VȪ�sZ7�ҽ�B��N�8ߡV1��`�F��a��DSL07ۥ><��ژ�u3�-Jce9�N͖(ۍ4ֻ�h�ߕ4Myؓ�@�_+y(���kJ�����/��1�ij��J��g;㙌���W��v� 	f��Q�>{�L�2�����e�t}�q���c���UGZ������~T�� �5=-�R[�v}j�>��ք�Uvߓ�͂�'ӆԈ>����?���2
,Р'G-�-�lRQ�B����
N�!��HA��ܽ���(W�0:	���"�����PU ^��T��5�p ͋2�^zV�8J��b�X�m�U�ve��^0� ������6������,��"�H���a6��c�!}��u�
�
C�BU:R8?�?{?��0a1� �[��п�,Iկ����`��͟@�E�/�փ�0����vO��������վ�b5���O�y��X���EŦ��x��oī��"�Y�Y�h�m����	�p�2we�L�&U��Q�Ɛ�ZZygj&�r~<���:�OE%A�3�s)/�����֚~���|;�GD��D�{���V~�x�C�Qc�X��G\��!w��@�Y��/�a�֌w���/�ʹ��#��b�yY�1�]?��GYp�ǽ���h�D����/��H� �2;*��{��b�G��j��6������&��o"�>���A?ϛ4�N����	���1��Q�����b�2���UK	G�^NaW��ؿ*
f�mp�(�1�\�����'E�\M-?��˲��b��<8�8��}�!<w�gN�v�E��ir���IҸu_���ז�lVj@ŀ��<Եjc�3$�ǃM�'ecM��a.rD
�έ�y�GF18Хta:d-S�!�̆��+����_���;�D��a����e$�'��-SP�)gR�u_��R�*�O��b��8k�~��NLq�f��G�(b�;5 d���.
��S�Bi�뻂� �� ��O	m�d3SN�[ظx��ý�G3
��tY����:�l���@���1�����<]Μȇ�=~9\IT)2��`>�eV誄�v~�#�Ru��
�A�}8���P�-MK�_��@�.ͩm�����7�Ðb�FZ�~.�k5@/%�v6o�omН���������GΨ��!,���3f
{N�v��-�^JBP��5r>��F���(�BGY�d˛�]���$T8�GK��+�E��յ�#`��
�*k�1��1�Ih�
] ���I�N��VD/G���]L˦�$s��b�X���D���#I�|�'��+򋎰�%e\3(�TGq(��睲�4����t��x*S���Ir_�"'���8� ЇJH���{R��B5�ω�0/8'�$LV��S9�������Q<]l»��ڄ�������goq����"D`^�\`�1����!�+w���J�+؏�[����T"G�
g�F��}���2JTC�~����|u��+��9�?����+W0䂩K��J»OL�
=;����I�L�XؑZ"9�L��a?�#s�!�U\�8�6s<��<ӊ�樻0+C�Œ��H��L�#9��wnE�4�l��Fځ=�1cT�s�7����'r�!am���
�?i���C����qԊ:YDI^'m8`�҉��4e�� ��s~��&(�O��՞��&p��R�uiV�[H�5��(ߝO,��'�|�!��nKNFs�2?1#����������O��UD�
��~g�0�� ����J�|0�-v����kC�z2l��2Ɇo��䲜�%���g"�K����%}*�`�M����ۡWb	�o�9yZ���o�S�����m�Ӭ���iH�����h�S�����^T��%�;�É���TO1�S9q�����4�J�[�A�k��!S��ϲ�&t[�`���}�d��s�Yj'�y�]�� ��N=��s�]��n��υ
���_\�bŘb�t��$�σ)�������vs���!B�[v��P�R�4����WF"��L�D��c��
�v���4_�d_�s(\�[�M����UP�LXp\�?��r]9A�s�x��׵~��^����@ύ6.R�&����B�w�iý�+0'cŲ?6�O�S"s;d^�GUm�}9�0ݜ`���/�i8<aT ����m�\�5i����C����L�r�AO�M��m�%���zE/G8Y���A�w$���q��ZvNQ�8�9P�jP*J�}T��	[j�� d6̪xK����H��������#��Fj�H���$�J�K4�q큙�;@���`����k=K7A������F'༂�������.n���y�ĺj�\V̷�T4�U�vC0�h���I1�L��+iE�8���������A�Xw�G6f��f��r�� K��LG�
�9��'q��Sw;8��k��L?�$R��:�b����2V�(4l<ޟ0�P�S>kt"�f�l6�QTh�&WX4Dq ��87�Xa������J�����C`+�J���õ8��lTebJoX�ٜ��f��v5i������!��Ė5�=N��y~$�Evh��_�6�Ɇ�J�+=UG�/�-6"�*+Ü��?��@��n�ܳ����	H$��g3�v?����VS�B�)�9͞F�l~������j�������z-���4�B���b~½��.��r`#XцZ���j^�T.�UZ�.�S�?�w˒��(/ %��[����&HEĘ^BT@{�2Jý]��6r0�T��݊��e�4�J ��S�_��M���UOk�+�\�Q-�%)�f[ ҭZ�H+��H�w��Tp5�٥l�+㏚��\ewgշ��X�z����
�+=���n"�o��^�PȮ~Be�7�,u���Tq(�-TN`���<G�҉��V����?%Z��'��>D�K:.�J!��%֏���!9։*Ŋ�K����X���Ǩ3!!4M��݆}18�֍w�`	���߳/3�SJ~����$V#$�$���@Sΰ*��a��0@k�h`�I�'*v�[N�iA�T��W��-���\�!7�9� W�
X
-L��1'�� 8��E���+�S
BcR���p[���C����V�JN��&/)�(�L�TQ�m�6=bX��"���i��n2#���Ƃ��"��ͨ�����	_��q��U�t�㹤�.�4g?��xf_���U��z%�r�k�,��_�w|��!q�� �����Р��JvwKp	���E�k�?����^zE ��� ��*���k�S/��QO"HB2�EaS�q��^tŉY�>�ǂ]��Q����qc/�+��{����*b�Z�.�;�d��#Hm	�d"�c��f���?}�*�e���M���f�Cǅ� i�Է��Q��/S�o��@�?]��k�'"q��d�*�^���h�6���;���p9�X�5��N�>P���*x��C>3G��Jx4�ޥ���9�,3{C���_�'�'�������(#km�ͧU%#ujZGȖoc��5��;�1����	�~�ƢI���0�upsذ�MP<ȗ<n��֤��Q��;��y�o�/V_��!$�7�+K@}��[�SX��8�<p�bY�mE���ɍ,LƜ���4�\����y\ x�O�c->��=7��[�9
����pEm�N0��E��ߒ��� >"+�����Oe>~mː��Y��N\#���m���1� 8��<0�hG3[%V�@����R�b�rӊ���sH-*�𔙥k6�s	)jp�� �$�ZZ���_R/���N��p�`���������|� 	u:Kɂ��uA�{��f�>~P5��eZx�57�a���a�ey����s�V�&�����s�C�P��vٿ@��.h���H����T�����@�R�l���b`uۻ��-*cfh�	�RT��zp[8ϸR�!�2�tQ�_q�J�܃C�zT����֕.��hJ���LR���	��S��,f�t!��%&{�$���#�S��-ߴ %��$�Aί�Ü�mP��<ώ��3L��3�����o�}Gi�c�K��Uc8���`A�7��fY��ÞX=�m�ֈ+�)X������,YHȼ��[R�N�b��X$}N�V
�P�����`%<���f��j�@���~�������	��S���������(h"4�� ��Y��2�y"�>�C�"yUCo�1�<�d��%�#@���=+�X\��!uR��ɣ隽O�e��#��䤲�e�e��ȴvM��s�?_�?����3��Ȳ�wk���M��\�2�ԧ��xMz�,_�'�x,�<����Pu?<Q���N2937�I�.533	
FB�T�MQ`~�_nj�F�պþ�����8B���`��G�a��`�z��u��u4�@�aꁗ�.{7+o��u
w��E��B�k=�@fZb�s�~�!�
�;i�^���>�f.W�QE	��b�r���=��DEf'ν��b������ꁺ���n|��j�7�<(�
wXSn޹V%�7X�Z�C�Y�GM>'�ŋ��E�-�UUh5&����$V����rn*�|�o�V�!5�%������E��l�KW�e�j.X�kR��x�����(ֲ����ơ�7���C�nZ`B.;ѥ0������̪��+��\�����Od ��	��� �O+N}w����T詄|���]w;�|%���nlz*���8=�R�ce�Y���|켕r��w���y1rY ���{��B�q��*��t┧�{|�eK�(��n�8n�
@	4�5�� f��� >�Z !�w1�L�Kd�ƃ�%�P�i�s�K�>�P3i���#]�W�E}r2	Fs�N;�?��z���9:H��PqM�	GLeE�!j ͩ�����+��GD4X�R�K� ���U��7�x~?��]�13��g�{0X��I$T\?��<�	���=6���G�t'>>ZK�+� �6�p&�
�q9�P���9����5��^�Ow_7�zRE@���O����7#]M��R�!82�U�����N��L�^�eY~K����z7Q�W�@ԺP��H�{�!	��]�0�Ë+���6������O܉ԭ`�߸+��^�J�"�օ#h�54�kJ	�ޣ�i����ģ�W*��L9u�a�� ���>�d��He�����n^���оrH�缛���XHg�̿ޅ����v�/��N�\0k�2i,�P�g4x��m(v��L�ј�w���&W����	������BF���TۆVi��x�>}i^v!�{��Pķ��Ku���Hv�� ���iǊ��w`Wʘ0
0�";�D2�=��u�k��kA�Z�;��U^����VV�1:t��]���m2��y&���:��4/�Ng`?�x��Cڏ��N������T�I'5rE1,�1Шz^	�x{�j���_��\h��a NnW�0�A�H��=W�@&�	q�񔬏s�h��6N,D���)ėjZj�@v�k�m�P��^�$����&ӑ���A��'$�Η>Ž���Q�G�ڟb]�&��H©s��l���t��k{\&D��Y�W���W�9��:��tP�2Բp=�(�[YK�-�K4C�=V+U;���R�`�Wy�8�̓`1~"�
����"U[�p����ᶌ�8�=|� g�z����ԩ�]���0 ќ2���Ү��"�JK�8��e1B�}z��>��5�UG�D(9!ݬ��"��Z\u4������:��L�D!G	��	�m�T�S���4
��O�%5Lϔ*��ts,'st|Zhs����K�ЍUl;>�: �rI�!���S�Zۗ&����fХK��Ͱ_��W��J���rG.�=w�nz^��m�ց�����F��i���0��G��Х��kNH����NB�+_u�ɼ��dZIm!`h�ġ�P�4�| 4Q#��J�e<8��إ����$q��Q��O�S�a�FD�d������S��m����
���RD�F�.q�o5&��'��۰�:L��
o���&�����v0��md���%�&�sV~�E������x?Ξٔ�h���	����k׀�(�L�ߤ�ԅ�q����q�z�#�D QU.b&�����Ռ��
����\�o<��	���U�����)>~��?-�^�.JVR�8N�$V���`�Wpj���GҠ�;gN�;P5�'��ɡԮ�~��u�
,�Bs���.��a��w+X&���R_9ȵѰ�#�/�V��E��}�=����s�a/ ��Ԓ�����,�N��g� �r��Z�(�_��3��QϊϿ$��6��"�/~�%�?Lp�������{v��P�='�#Ј2�h�W��!����$���uO�,�%��'��/	����Y4 ���G X��ob��+}"�ή@�"s���rM�xi��������H`�|kG��;~�q����3�^��	�Ó�Xv��q68��,�g��F�+yD�Nj�`���!�Ȟ�E���ϓ̺D�`x��՜� .+��T��A8(�kl�.��f��V��nu���Mhvb��@ުl-�b�܈��L��Z������	��9'�&U�^R.��F��2���;#�Hn�A�k��G�/�g��v(
Gb�P���p����?8�.j�[���&�Y�#��E����P�T��h�y±U��B�w�D�a�%`��8B�mN����z��Y@A*�����R�0uH:nj�,N�"ը�%y`�����.2��n��.��Ψ6���*h��:,v ev���5��Vyu����[�i��S�_�xޥ��5�f$ <��(��lFm8EE��7�ذuŧ���L_�]^ O��߄��K<�n�K2w*��g���*�S���(�n�"0w���ZI� �E�~�=�'��>R�V���BMO�l"��=�V`v��)�3��Y����P�X�L@��}1}e�vEY��ع|Џ]ZΞ�.�	S�epg���_�1�G1��(��dj'�uu��g;Xۆ����)��sB5�J�a.���*�s�<�i=���k�*8��g�V#/"dQ���I�K-Gjny�sI� V����i����<�����
w����L����W�7	t���߶uB_3u^a�@�!���D|9�G���$�F���%
[��M;%��sypS����e׈�a@�ͤ�� ^ߺ�2�U{�	����pU�QT#�l�*��wf%�*�����ynl���Y�� 6�͋[�%ѯ��W�9��m��;�6ڎ�	i����.�z��	�$��\���l�������X1nY�lE�B�n֎[����%5Yƽ5�y�pμ��pC��眽��9����L��C��n���_!��6�᭝���n�		�� [^\]y׶u�9�2������Rr�-�P���Q����P����!d��*k�ȡ���z)�8MR����¾_�%G��b����s�A��'�"��ڪ�W��u۷�?TKM��Ӯ`nٗ&l����@�[�o�L�����G5y�]���<}��ˠ�Oᩁ6\���|���u��ƃNڎe� /��S�<���u�c�.�<[���*��F�@r�Q�{�ll0�i��Թz',z����US���*S
x���[���S��L{�
��m9: �c���5�ڿ<��+�%���<n�M�`��Y �aǿ�?�����~�'����r���Q�*v���?6O�^�{��/I;]>y�����+�У̹�����z�Ve��B^MĴoNv�WԼ������])P�'�Q�l���o�k�3�-um� ��k�J}:|C�9	Qp;��k��D�f�֊c�����H�D�d���YiB�0ϼ:�ȼ�㜛G`��p���x��.�{x�@Spf1 2Y�Ҫ*����H��р,0�%e6Øb���V��I+EC�UmWK���m�R#�3g�Y�jL���j^b��Aw�G5�l�bLW��Ш���;���5���$���4D�J��M�yF/���s.o}���?���3�@q�Av��l�z�x2k�UiZ�4�D���UL� �[���*�G[8L�8���	 -t�������J��Y� �]7z^8_���1��B䠵[<���Lb�$X�s���$�4� ����ߓ�O�s�R�8t��sP��?�[}|^Rx��1M��Ꜳ����Y[�$�0U[�=4���R��-�}lQ�i1�r�lˬK��kit�V��Sͫ�u���j[��Jޙ�&�9��y�%�H�G/��8�J��̂��ƥ�鄢E�fH�E'��R��6DL�o�4��+��U�CÞ�r�4���D e��*�i�s�bS�zϊ�������zj�1���U!C���>�d��j���:_X-D�c!후;N�-�d���0Ђ~�8�����eV�.�L8�D��+�'/46�lW6���=����\�T�ϔXxA�T%����?i�19����K�_9~��PEU-4བྷ�+b��}ڰ�.�� iT�T�G\y������n��I�H����t��}�/�xF�yo�ţ�,�zN#�l��؜l�x1sڕD"�
9u\�1��=�����W��z�KH��)N�Qd�v�I}�& ��(���g���iJ����(��,��E,� v��9���9�ΐ���m	���#��6�\����)�dk	?z��>N�ä�nڇf7��:��ɎS@�r��eo�!�h��lm�<a�#�u�Ŭ�	��Vܥ#�̍�{��R6��^����D�V�6�J�ő�(��Ŕϵ�X�:��z<���Qk/jYx���ž1_�U�E�J�9���M$��ة�!h�=���_-k�b�i"X�x�sx5T�0w���A�0��E{x+��
d��2����+�=�n�i4?��o�l�T��&tmҝ�~}`��R\�S�qx�Щ��@���ٯ�����'�����@>٘s�0y��ˡ��+���Y��~#��?Ҡ�#a�+�t��3�5�Aˈy��-瀖�����7W��RQ -w>��.�R���|�h"D�h���3�7��dK (˘a-���0F?Va�>9xQ�8C5�d��[ٝ��*�L ��d"��x^g�֦/8�m�>P�Ww���>�/@Ӌi��	Fh��}1���1��e�tIl��hBg�ߌA7����ޝ<6C�ȏ�C��:Pu.P��T��)p�gtO��8Y�S��9?0d��E��q`i-l*�<�)yjX�i�8���]� �M�P��]��~ȶ[�(��2�m�(3,�p��k;�����BALVr� ���:=�$�x�q��j��ڮ�z��9&����i�"78�5��$s,oCa���?���+�+�q1=20bq�ddr�+��{����}�e4�K����M�r��d�,���H�2]3�ߺ�3n�fF�҉g�5lO� ��c����ʠCR�$��py��h�-�64"ul;� ���eg���&���r3fx"�@Ll�E#.@T�2�247C]�Oג���忈�K6��V0�F����x,�t��a��W�nl�Z�技S�VF��ȅ��x��b��`��V��2I�Q��K�"����¿}�Q�/� � caF5�����XXn�_/Ť	K�(� ��n26dl��'}Z֥�-�g_�]��Vʾ��e{|��Gy��b���I�=��Ɇڳ�k~����D�=E��g�V���tI$����t�@�uƫg�8��i����tx��� +]G��/��YsDNr�a�a~�?p?�7���*$�kd1%Y%h�m�_VZ4��%^{[���/���
��#�8B�wJ[�Y<�\���i��X��)�L_y߳:�f8野��^o�_�o2�MgU�^1 �R�9׼42X�A��91�R�"���N�������{�Vs���[(��/!wq�A�ڧ�!��Z�e��uMU��:�rkꭙ�+��p0"�UHסY�vQm��NP_>�\^=xw��1���_�4���zZC�>� ��b���/G��}6 wawD�N6i6�Xc���'\�c6"`Y|i�[r{���SZ�����|ѐB�)����-	�e�YΘ;'����9
���s�߾���
��;gTVf
�p�3}��[C=#�Y�'U�䒖�hz�9��d;S��xڂ���x�%� �����t��Üݷ�����Z@6m�����-}~��0�*t6�~z��<si�Ԗݔ!��Q-�W,_+O9�2�^f+X��HKb���xH0l�3SlM�T/;	�zF�~?�]n%CE��0T]_�-f�A�/�Z�wgH�7B q�<k�AY�GՉ��=KC�DD�-��[�5"�O2�����3���Pl� ,��J$u(N|0�t� ���zԞ�&��ӤN��d����in���\�]�֡@+k�֙��T�-8^>s��R�ރ��z�Ԁ@���`�2�,g6�>� ����Y>7+��Ql�G�[ހ�< �6`�/�
��ߌ��W�M����D�nC)(�HhP �o�a��1���GѿHɕ��*�ĢEs���G4��M�йD��r�Ș<p1uaV9���p��$LXR���1�4l!LB�\8?i��ޅ�c�x0:���)�������36���?�U���2>&2ꬶ��t��WM�\`M�?s~����
ײ3<������/�Չ �=�� KO�-:��2�'��&�V�6�35,��n%�䙧�G��w� ���D���$�g��o�SG��ܺ��I�ͮ�I�ƿ�Ba.>�3�����@���qPAX����	���	�:l���U�",�˙˹i1<�������6��������)��-���j�H�T����UN,JOCӆ|$�
%z�����S�X��ʪy��,Hy�>��{RM����F�  �N�V^���Y� ��Јðө	�����9 6a���qF�8wl��4I�*)�"-�J����3�ِ
ñ��N�y)�aO��h�.[�e�"�����]G&�m�LD�L�^�V�R��K��f��S&b�L��{�83�0�����\�w�_���wvOw���K�n��@�������Y���f�^d���g��V@�OW��-|���T\e>�	S(���S��[�Ӹ94}���O���6�.7vkF
I�� \A�_�	�^_'m�Q��U5OY�7*L
��%�߁8=G�A_�n6�֝�F��,�*9���鉌k_�t0Yg��-��O\P��)����Y4�Kk�Ǘn ���ϛ��B锾ѓk㗪�Y�Z���X3��M�X��ӮlE���V�ޙ~��o��r��
�˜���_��	Rxp-�q}3U3ɚ���(�lL-�~�D%��s��v!!��3hއ�^��B���_J���:�fT��e5�����oO��e�h~W�R�;���&~�I�g�)���4�Y��A ����#KG�}�/�W������^x?��JP�0 ��qs �ʡ�阬�!�����0\�R�|M�
s!�ec׸{�c�a�e��5?i���;fS�c�1�,Z! ^U��6���cn�M�~l���n�q��a��ᣣ�\��A���Og���4��4���eO�6�1��24)�e�߼��.�@�P�ܥ���+ʜ!�|	:��P/'�)Ј%D��6�K�&< q3����A���9V�]C�o�@=m2��q� y���4a>Ǎ ��{�W����V���Jl�f��z��X�
�7�e���8�����r�Q�DW���������SP{��Z���c�����E�;�F²C�JOmP�$=m߈'��A��RA+=�y�@k�7F�����WρS�8���G���!������l�M�D��1�Y!�*��Ď�|�'�.���kMڸ�����S�f[�)�!.��wĭ3$B�uM�t����8K�/�D��EAD������3�r���ŝ��b���8�:�[@1�/b܍�p�P��= gwExh�[�qw��Eoh�s��d���(��Դ����	�XNQ�5!)p���'���\��S�*�߯��{���z�ŕ9�~$��dU�ϫm��f��t^נ����� �7q�Ѡ�%{X6��T �,��ɘ�		��������}H⛠X	Y)�37�e;|��,3I�t���D�E4��� ����`��s�j��Vҝ%+��)�B�x[�z{	<���)������p��獰�D�*O�h�ó�`
�MF�>I�G���5p�8+9��v�k�	�,���s88֎�>��@���p�@Ԣ����`Ɯ0���t�`$���h���6�-�+�5aK��}nҥ��vg�}�3�v�����r�<,OWi�T���*�8���ī����#�A�u�3<�ܗK+�_�O?�5dkh�pl�ޠ'���A#���Ub;�5
xw����窑��p���
iM�h��G� 5@S{_��� -,���+��-�E�qgYl7�FT��B�����"R��(�܂�l���0��&�n�%F�Uۃ���`o O�K[�������K0��>�Ӎ:�/�`0����|��;_���.ɪ��R��8Hi��Cˇ���~\�.K�P����wx��2�b���FH���l@쵧}� �1�\��/없�&h� �W���йD��K��Ǟ^z&���"jIÃ����?�_<�Y�J*�kZ���O�����X������+��yk�]�����އ��ý1agL�>qlݷC�tBE3�&L�;��,��(��G�~٣[�īp�����2�^��Ej���Z��sؕ�Y�<�6>Ӆ�гj�������Cϊ�M��c�p�����U���
lv!�W�t�iMHk>�^gM�@��̎Rf�E!՝�D�!j�]�Mh��~"���7�Gn��ZuQwrq��>�:S��%nkZ������<�	I���7,}��D���4Cj��C��}قM�MW$%�qx�x�`��p���B���&�� ���!NT�j�
����S�����I��ƍ��4��d��"����2�T��rY����lw�<�_�)�~[o�@��@��?�m��M�ژ�ډ��V�0��l!� -���f�^���=�� ��Ѽ�P����������u�2�kW7"���C�>�v%�}�r&��q8�^x{6ݰ-��'�[��Mܙ�n��I@���RR�Y���f�wD)wfw�A�D�,��� �#+sv��j���v8܀.yۣ���S!m9p@^M5+�E���n���!9����kv�H|Y�����5�B�Pc��L��Sy�v$Yc�dl4w4���_��k9��Z�"!A��%�8\��_����>�݂����>�̙2���p�l������QsLƺ�𾵆�����g���\#HÇн��1��ƃ���rf�Ę"�{х�	��7����'�k.� /F	�59#�NE��e���w@l�E�����
ʺ2+����!ث���{�}�f^?��a��b�h��B��tì5�a<��ҏ�x�1	x�|5aO�a�:�8jѵ���@	�˺ݱ��p<�BhpƐ8��VB���}G�� U'-$��g`JŜK�}2���x�f=8�[Gp�09ƖxV���hߓ���^�x���q+ͯsź���c��X��j޸=�����F�H�N��,����(!���/?� �R��V��Y�W.�d:
��4�xa��M�:�b�_.>�	tv�8h~s�Ki��m�����u��7`6q�=}�DbX�0k�ڢ},�\�6�0��ޘ������ig��Sj�#l���n�Ir�F���0�����ޮr��Wg&�� �^'�Yh�������u���(�Y�XJ�|V�̉D%v*� 7?�\W���=f�κ���w� �޴�Il�8.F�^2H�.3S��+��=!�Dk;6��q	^����d���q�A�}yR�*�@�.Y���b=>�՟H�>..e�]�)��:z�g�ѷ�Lz~o�
����d�
���������0]N`�'`B��46;���x����4�FPA�C:P���e\�oi�3~���j�9ϦO��c���8�;�M��G��&7��Z�O����YCun�t�23׽j�B4ҙa0�1e�'%��aފ��e��g7��{IJmIY�޹$�c׋8��{���b�	�H�_w�3����W�Pbl����!f��G���a���ꐹ2���v��\��5B���^me�Dio�R�D����\�<`y3��ͭ�}G�|q!�x!񍮴���4�gbG�ls6I�A��K��5��?����x�Y�wzk�;c0��$b��+�$�:��yo�Y*]$K�Jz��v60��t�g�ף��x;��g0��i����3��������]<�6�]Im�z1ӵ$����c,/&�1����l�B�ޓh�T��T�琬��29i�z��ԑ�V&7��DW/�B��-z��=Jr�1"��-�&�3C������j~�7�"@���� #q���֌Es��bxmʢKZ�S�+;˗�9}����E5�Ph*/�{�R��{����,^�"ic>�z��odv|�;@mDQ	����z{jo�'�G 8ɍ�wb.$����-ے24[�Te�0�a;�	���ZaH�zti�=��8+5�+�Ċz���^��H��C�%4X��ݿ�1y�z����i�H!�bY�a���X����𢠤�b'�m�[tG8�Њ�l��k(Ib���~ʼ�����oV]�U�luU�<��]�
5�W7 d2'���@\���R?Ed̉Fޞ���!n�;iy��(�8�MdL>�.�S���{��0�I@7�߷"P����]��۟�A�j�3a9B�p	!�-���ծ,H�O"�5�\�Sd��~�-;�N�dqq�2 �"�U|��g��s<9��NK�ʶ9A������ MGz��d�|�=$`߿��b�ʑ H[�UiU.��,�#��������7�0�}�}��҅g6ս���C����iǴ���u m��~��qo�^
y3���1
����m'�>d~g�ֿ�\-VkqR� 0�z���x�88%R����w���C�m��8>�0?��O�ٖ�2����{i��U�<�Y>i���]wC�	P�zĬ�����1)�O��4` mܦۈe��5�l��$�5)��ϕ	�5�N ��M9����z�dc�ĥ<�}�F�O�y���ٖ���ZX��)綊 �W�6/[Vh�!�s2�cH��p~�!N?@)qN��������>���I[~�{{�m����֚v�Whw�5YUa�)��� ����h>9Jlx4�Ǩi'��E�t�	&�ێ�]S1{��K�ɽ��"��Dr��C�|�!]D������
�2�~�s��ƸU@�8�4��#�t3��� (�G0���ʩY����Q�)�$�bڢf �r&�!oԚ��R0�D�w�]�CΜ,E����^��Zz��5Vf)��pX��E>׎N����*��0P9�Y��e&9-��G 9��-3e�K�b�i��ȑ`Z)�(L�|yH椞i��2p��8f��!]�G��E��O���OLl�z�U�j����0�,D�~�b��#M>x�SLeeo^R8*�*��0���v[H�"��~���,��t����Q��$� >-'�a��Q;�g���O�eD 7���d@�7f��?���l5���x�'m�k�}��+�����|u`�� JZ7�Ƅ�R��
����9@�t;�`a�hN����v��x��=�N�[��H�ӕ��V���Btԏp^�51�'�o�I���@��^���CM%\Ξ�f�i]�|��6湒��fF��0��^g�hr��U��������m��Pv�d�α�*�rw'�%�u�G�}�ڟ�b���D��n9�f��^�2w�/A�,�&�������	��#lz�u��gUt4�c{x[�=�i	�r$�!�Y�2F� yc����8�߮��(�"s'MoB��@��u���[�`�A5Vȗ���/2d����T�s��LO6?�.�0ØqPqN��-6;&�܍#3G�uB[�DkV0^L)C��x@J`��1kh��H_]��4�d��0�d:A~Z�'b~2��S���V��XH�A�L��Ү��4��pwyg�^/�[���+�l|�{��౪p�
��:�!"�����vv�"рf�ql���D>����vx�é�ۃ�ۯ�Lob�%��cnhL��c�A�}JkHm[����¼��kv���3	n�%�65U�`[��I�b��!k���6lO�5�v��G^��g�F�<�c�Wc7^���ۄe�������_��ڃ�fz��� �fA�+��C�@Y�9;nd&�q�{y���9�lJ�Z���{L�Ƿ_1��+f��؛�D�=�<O�A�R^|��2&t@��.^�j�v�خ?^��`��f������\eU�$t��햧z(����Ǟ�8lGt��j�8�������R��	CP��G��I6�3�}u�C�h:E��.��y�$�(g�~���B���ac�A,�z�,�~��/�M�Ԋ;�-���j��Irr�aG�q�U)�IF��'�=��pz�m�������\h'�D�]3��M�%��QX��H�b�H<&CH�����J����#���o)9<��wN��m�v��9I��U��vEv�6 @IA�2���}O?pT3v1�c�k���9�wӤ�������me���G�6�
3��/�'t��]�L��Q���ʼB�%x,����Z�-cH}�C�����a��y�������Ұ�b|�YK`�4%4�:&��SD00B�+ܢ��H����p1�h5�ދdn�{k����%m��C�;#ĺh�I��<=��z�3�p�ʌF�L���X'�R7�������,&�����O�5Q�x����$}1��)��g_#y�c��U+Z�-��$���A�>���ϑ'I�v>p�L#�d��N�x��#6�m"I�����:B��5��y�k�~�1Z"���[(_��W�����Mܜ3C#S��.hK<��_�������<�KNS�w�~y������*�A^���	J�＊�qi�тs�*vH�3�������Sj�s;|����t7%�ՙ��j���k�<�Oi���M�l��8!����]�3	>����pX)�+oRO�1�Cm��Y��"F����wK��8��1����v��g�K���0c1����H���1�i����-���<��i�63��� >��lX�D�v�B9%�5��֫������4�������ש�L&�;2w�Vi#d��9��F�8X��>�'g��ʲY����Ne0SD�2̡�;@��g�M����>5��R���D4Z�G~i��>
�I ��[�?=a��E�1�dop���MA���V��1[�#
7��x�������%�`�	�`1�u�x�l��<���@(�!uC�,�z��<�D�a���@2�w�ٕ~��h�nrv��p�5l��T�5��=W]��.I���Dk��D	47�����iy<�������o���,}s��j{&n�\j����D| 	}*�a5�į��q~��/��;�Zj���i� <P���,^o��$z� �[{�1�,	t�t�q�Vq�E13�Y�qg�}��u���y#�z��{��?{y#~�*5M�d]����ߘj
�e
�A����T���i��
���O�01�R�o����̚��$�Ъ��@�6���,��v��f�:\��A��`�W\�VD㯨w�qd�%PQ�A���2pB�?~h�$��PZ�{D�t�g4�*�n�`�-�
 ���yJ�%+���`�)tAz���J__Wak�ͨ'�Үےl��I�h���s�}n.�o�Q����'�>�����
��=w�^Ŗ4f�s������ H�o��\Zِ�f$)�	���`��b�W<W�?B[\k��~3��6���!ZBSB����Z�W��'2�2{����/yBUZ=G�wq����-o ��_�I����x�E(ؼ�N�ۻ$�_�\K�F����Z��"���vU`�90��6�h��`��V=@1�B�u#5�~�6����d�8�:��O���Mu���#+*D ��B�j�M��u;����|�J���^a��Yt7Uق"��#a`;�(SP��A��U��V��&�*��4�kܜЌ�,�y�����/�� �TI^�<����j�j8Y�y��p0���O��$>��Q̝qA�����ʚ���uA���ѥ0�]W�O�Z=I����To��ݡϮӍ��R8���V=�v[J�/�:���R!��>/+� �	�T9&�\�9��bbT�o�QV��$hU�唻'�^j���i?�_�Q�\���k֯�cM���%\C�сܦ��.��Ȉ�҆�m|�g�G�q�|P�Vr�'��q��Zֲ-)"vN\2�@��ϟ�����%{�^R��M7J��xz��ds)?Њ˼��)rOI/Q�2�a�D��[��ۚ�S��]��͉�2\]R`����(�;��c��֋ �����L`j?�B��&�x5ZU��а����}����ba��;�{��b��₎߃�f�� ���q>`-�N*)�>ʈЂ�e&`�3��O`޾��A磾(>�⺲��L�^���� �@��|j� �,{�x�2�V1��Ƥ�&�H2��C�g�շ\E����nc��3�/��R�6�xY��K��黭�.��E�M�$�|*�r_�g�w���f�=��;��_��s���)��<�Ϗ&���/&dPgc�$F�3��՟w@�'����F��cv=������v=A
��K�(����tGdZ3a�*,(�M�}�i�Y	�s�����'�����I����3��\yώ�[Y`�L��u��cW�'x�$�[�$OO��'C�qt{�v S-E��K�s���:Y��
^]�VK��C�a���S�Q���dwu�3rr?��V�2���b��}�O�}N|L�_	�u��<)�-zEi#,h���Mmסt���IS�W�)��������3����;{V}e|��� ��\5NJ���x��B4���p��8c��y���|_���G�Ub����y�سk�m�e*"���7N�+�q����i�4iYu8�ոE�t�ߴ�r�NX�ab0�hq+z?X�?�#�%J�6f��\�(��̛N�ˑ�6�'�k��s��s"ʜ�x�����F�)�f2�n�E�u.���QG�M.�s�eR��L��(��Q���,�p
������>9�#����L�� ��c���S��F~���Dz*?z��@���x����� �־�zv�Lr�w$F&3�+3R���w$�`����&w�dy�#s��"D?4]fQB�����h�J/�*���]�%��?�~���K��殞ʰ�����H�;�^)��'���F�7@�`���������Vǎ�q×�mR�5��ֵFft=C�a� �4���E�}��wl�5r�p��1G�����q@Y���7d]��;{��8�k��l	���̒�HQ5�� %H�������H�������	� %N��X[ ��[$�1�g�U�����F��?Ǥn�����iP�jX.��|�+s�D�a���(ɊA_g�G����Kc�G��wF�x� $%<9�J��M)È3C�v��UM��0����ڎ���jۻ����� ���jZ|��ћ�Y�9l�c.�E��-rZ�3�̶E�~�H�β��/��$�2=�+67���3�"�HC��f��0����TKG?4��d:�6���S�Q��� 9l����A����3лU0��Ԕk���.kU��3|Tb	���x�N/��8��t^��?���)l5����.��)��r�[j�X�㠢��E[��%�º�@�}&��!���� mo�po��D�!�j�GKyH�|JKڳT �v�MTh%k!���b���ئ� �Wr�uR�;�%M��\��U���l�=�QZ�A	��Uk8)����L�rX��׃�0;jqp��&#��͟�ʧ'P1)K0��s�=#b�.�:�1t��[(��P�
VȦojV)s9'�~��V]ԁ}(�EAAN�4'�!v�4���:�~����sD���"���y��1ql.���l�V�R�y�]�цH�Ze��9�k�O�֮ƣ601�w�Ԭ	����7�����?�Aw�q#a�A9~�}�,��$��D�8L"�Ca�GP�D!_��g��wI�,�~5�v�e���������ɕ�<kx4�ÖJ�G�;Ht�$߉E�~�;��<r
l[���F���K9���C�:��� �eC��[_.e��Wƅ.cd���.O�9
~ui��$�m��ɠp�W:�J�,.�|\�T�����U�S���I�6a���DD�pp�Mib��R��k�4��`��d�d� f*i��Ȅ�O�O#x��<��Hhɶ}�`���Xh�gV0y�3Ƴܜ��hj_��ǹ�;QAxx�ଋH���+_�zq�i���9�$��;� ����)sS����{��-�����@�[�T?Ϙf0��m��M/ӈ#�k;���//Lb� u���L������6�].`11����&��R+�&��Gd��(˗�k��(����-Q��V�oп���߂3�Z����)�@&�v6t�q[���6�T��]�(�Lh�D��p]�b���(��a�ȶ�;ٍڶ�aGIXߐ�!h��t�^�s,����Ȩ� �x���={	33�i��@�Oޣ�J��`��j'#"ݺ����eYW6�7��m�~P��DU�K���G��l�Q�.>�:q�N���
��̙l��4�W���D��MB��ŧ�r.��bʃ�{A��=�Z��w�1�ϮJ ��A�0��M3�E�J3�$_>ЀV�~f���k����t�`η���a$M�R1��Lw�+(
���[Ú��Z(�c/����o	���%!x�	ͯ����5�E`.w����q�;���M/�$�#B}{p�
�U���z�(�����>q�I����gn�6p'u�e�|���p�4r؅s%49�]tkc��N�,^c4^�/�o��F0`�&O�`Ib�FR���t�F���;"c���C�Y-�.[S����J^j���!|�aB�(��+���-�����x4������B��9/5�^5��A�LhI/�	�;�@T������X{f���4^��]� �Ì�K�|{>��+x��8��!�������	8pS�QJ'rV<�?����@o��6���
����Ȃ�l���6E&TZk��Lm�� [��]��
��IJ�����&q�����K�=��n�˿
�ӛ��<6�=��F� �
pf��E!���ZY�@)���{��`̰F5ʡ���t��r�	*���<ǟ��b�!��op�}{Q`��k`�R����|v~l�������jU��#�����w��� ��2����Q�{��c�{s(�� ���AvD�(��s 5����mCPG���3���*W�O�ub�!�S6gH�K�c���{ڋ�4/]�� 8�s�X�ͭlg�=������|]�[	��պ�
m5��t�33��.G��y�te�{v(� �}�G���:����t|iҎ�1Cp���4v� ��i���	wvv��4�V��^�O#�~T�����6���I��xK��;�Rs��	R���%�v�&�ᥐD�g��.s�6�ʜ��U���t��ӎ�ә<�R��
�7�a��J텧��Ϲ҅��|��`hI����a{��Y��gSR���x:rm�����������"pV��J� ������5ʝ[���q-��X����D�A�T"\�+֬�|��ܡ��}�`A�T[����J����B��<O�ZΘ �K���(���D������rC��6 B��䍱g��u8���ӳ%�^Y5�Z[�E�)|���Rk�m'T���\�s�x:1�n.|ևI��m� ������>�@�����	Fhd�J����9���W��&�BZ��$�hJdԁѼ�B��t�mc���nG;x�M��J�ň��wД5�
���;�D$��M�k���n^L����3��U� ���w�r�oͣ�/Ք�*'k�!CW�j4���&�j����;��!���b\2E��Nt��D��Q��C'�i�f���A@_k��T c��+����(ʬ1���4
��V}y�{��C�eN��x��#��)���M�Qu�EB����e�+ �G�]�>�uT���(��==te�Kx��#��d��37�_�'3�F������ Z�H퐥�!qTo~�2�I	�PbK�G@�FYڰ��z�Ia� f�э�6+�B-�����4�`��^X��	�Ӳ���8H��Vn�� 'Fu�j�id���r�g� Xj%t�����l6�&���_B��g��P�T&�u���"�Δ6�~�; zq�
����*F\3R�K!����{�Oi�"��dK�3zK3��MH��h;	L}
}�W�t���m�'x�р8G�h����*|���Xvu���g����"���8�p�O��b!)Y4)p����JHٻ_g|�fL_�fs���!z��Q�|39��m���_e��sH�a��dl����c���~�\�Ƹ-Bk[�@�9Ub����o���D[�^�h:$.4��q9����}B[���v��A���+E�f�>��n������M�ǣ��>oW��s��c�k`�z�)�G&�qfiR�9P�>�De�ak�S�k�ědz��F9h�X�O��	��}z̷�,~�_sq�^�L)!�ۊ"�K3HaP�w�W�r�efFW�M�����nl�,Ӟ˴�|t�����2+��W�sy`+�����vm� ^Ś`uyy���Jǋ���H*��3c�$�Ls#�V���y���W �?����D�����"�0A���]E�Lz�s���0��?@N�&Ὰ)�RK^S�|W�²D��õ��#�~��X�ó).r�Ƌ��+�j��P��7^䰄�9���⡐�Hr�(aG�fȭZ��^��b����v�ڞM�:����	��d�ІIz�ì�q'�u�}h�B	P�$�Y���} W>U(@>��'���;]�SX��[�w �o�ϰ ,�d�2����/ȳ!�FR�[.�s�	# ��I�^��¦��`��%�b�#��a��UɹOv��z�����,v�wrQx�fjӽ|��fR�gz;��'�@>�7]sE�q?�Ϸ���pmp��
("�Ѱ`w0i�kk�Me�2��B��'���q͟J�A*(���㛌W�f�?�����ܟ�JS��R���T�ACmAQ,�|N~"��q����	�}r!�#�v��k�-�w�ג+]��OQ;�;鑬GؔY�`ƒ�دd��N]4sB�5�C"�e�H��"<@y���Ϛ��j�U^Ӵ��=EUB骎�����Ev�2K����W�����+�S�,���>���R�[3�X>���X����ɊW�I�.�H,�9�bĸ����8.4V{���r͋aIʬ�ne;7#i�[�8l�M�
@2Ş�6ɔ�w|�C�)qC��~_"��nf��Q/���f�븛0ܵ��U�������<_����3I����)Hg��7����)`	��0 ���^���WƘ� �mkK�ic���p�3(1����y�+�*j�}n�:Bn���'�����H��"kX*pv?x5�^�T J�#��c�T����I���� {�53���Z�u�d84�Ls����G]��4��_Q�g5Zt��V�b�F<c_���Kq�U>�25x`�c�q�R�n
��?�no�����֡�.��nc	��<l�R���l����=�@�&a��NRځBW-��l?M�L� ,�]{���1"
��N��Q;="wd<�z��@��AF�V�v����ںMt8󆹄�W�����H�*?��V7I�����z+9^���pUA�ph�:�b�Wg_��ֹ&��$����0@Nv�@�8��	�)�Ps���O�G&5/?Σ��/�GG�T�'�%M80���W��O����yɒ$y���pz��@�"8(8��D�Z8���DB:�4?�a�T���c�0�+#/�h}��>�&t��#�OJ�Ua�CI&9��F��߅ T,�a �y�̐��4�#�G�ж����{x��t0�X��X\;�� �?�yTԁ ԊpU�KA���B �B�ӣR����u���%q62R�s�ؘ�gMџ��ɺ��d;���լg/vg��Y9q�%�9��>�ZdS�)��@m��o�v*#��?]�`����������b����:���I�"qQ�
�TwKY�tmţ��C@�*Rz��$B��5�7^�@�s��
��EZ��+����r�*�2��R��kx�`�gҹ�t�;�x�I��2U?L�����T�@���z��,*AR8�ì#)�A�C���~Rn��,�ˑu�Q����w�o��]2���u12�:޳�ʱ�g�.+��	Ό��>��:`�nG�J�ƅ�oZ�g5X&Qa�c�~��5�I�����SZL��G�c����Á�4dI-R2����|Ax�?-�Y��x)�6�H���B!�'���"<0J�y�����ot��{�Ǒ�e��<�N��h]���UM\���p'2�����?�n	C��)�"���.��8#Z�=�����>�E��}�'#r�� ���I��Ⱥ���?����B��Gυؓ��4�z��C]���~g �O蚎Z"a^�L_�f��q���Dx�TGpi�dt�r�ݸ�*	X� c���Ї�Ǉ�k4��/�(�e6A�r��Z"�݂:k�΂;a"�}�z���6]��~��saV'ī��;��<�+�K�!m� �+91>`��]�k1�O�ã�]S�k�a䂘�C{8��4��X ����Ŀm��a.1��@)�NOYK	�؃T .Rp�i��d���+YO<N9M���c�P���V!H5������N�d��4�L[O�w�p�,�>����y7ɸ�n���w��P눥0��s�\���w�����jW�
r_<��+�R���0�1�z����e��i*�8� �BMa
�
3\���K9�c��'t��p�1>��@T&/���Z�O��l��7�4��Q��X{s�46��"hfRщb�FD�0o�BRtt�<�����	�����e�Ԙ���c�/P�?�H�_,Nx+U� ��C��V�1��Ӊ�*�aax����a`bP 6�<�ҫ0�V��8<��Nh���	��>�%tm�}�+g��L�"0�q�@I�'~G"+ �	 ���.��䏓�<���2v� @���衍;�}��V�s��dHE�y�L*���뒢A��}��#�niX��*gE�L4���(���K=~?�E��*�/�E-�`1�e�͛�v@k����$F,�Hy�=(���b���0�����OHD
������E�����"8-T��Im�&�UoÓ@�xx����^tR�e�"�����iV��غ��k�j����B0�ݗ����_��8ՒU�}��e��P�9`#=�1���$�&_\�+��/S�����U��0X�m�h'i�&�d�Y�n��2���g9�qJIlW]�,fW��m����[�8|^a�����X�	�����x;n(���Wk�����J��l����m�K�l�i�T����s�K�4?ˈZ,�[d8NQ^��B�wPJG�w��(_�J��	�yFxpɹ�� ���C�:n�ut?B�z.�cx��r����RM��!�!��,�.%k�Sw��Ǵv��S��=s����E?�h�1x�K'�}9�����]����E���z^D,����.��o�I��ٔj��5�������(�.�5�o�Blj������0:����|r/1~o��[�ǽ	�p�-2&�ޱ�D����7�c�S96��r��n�H��s�_1L}�A�f +Gޟ��'�`>^�G���K�* x!�/[)(�,�&��(T�rYuj����f��d+^"��yi�,�yTw�~[
���[r00��8�	�	���I���W��{?:�2?�mt���'i�-�2_E�������X�Ȯ�|!A���p��S�}��B:��q�>� ��+"8��&�~��B"�PV�
�e{�k�1��`�i�)J�-���_�	���T�0��V㶣���l^4���W�<~"b�T/svi�c%�?�������ʐ_���y{���n"�+k�;%8��F�O�c2y�����bq�E��B)�p����W�*B'#=J���?Cs{�Yz�w���,�ɖ�I{T��ש�� ��FS�F="��*Po^[W=��˜ب�ϥ�� F>{�RݖԲ�'5&B�<&�
�w�����B	8�QR\�h@��R7���߯���L�����-Ǹo�O8���� �ek���52�[���~��*L��w E�Ȭs{�_�f�Qc����aRI��[��&7]���n���a�fȕ8_�+�й^��d��A�l��Rժ-��`c
�/�g! ^�԰h�ӤȇI��B=dҎ�S�b�趄�D�hv��5��/,�k�K/���+K�l?���������r��g�u�
�����7���ݐsZr� �jH;sp\�/]ܬ�SF5�W� i��=��a�ﰣ�Մs&�E-��)j��JD\�q�E���ϝN�
��?�;̰��	(h�@5^b�b!�_6����j�@E�0s.��>(G�}���l��j�57�����Fi���Ǒ�u*u, @������ّ��n�pI�A�)AA8�*ty���x]ȎE�ں<����s��O4��ǟ @�4�[�*z��H"U�B�~�{&I�����̤;d��ov��@W��C�^�!tqhs�r_�B�v�I/ndZ5�;f�V}�Qֵ�2���f={R�Ӑ_@��܌�D_�^��Q_�~k$�u�m��V������y�3i+��l��θ�z�s����!��w�_��U�D}��s�����Q�&'`0��%f�mk��Z̐��:�յ���8�TN�L�=��sͰ�$߁���=�đIh�-��LI3����K �=E�	w��ᘸ;����rz	ȩnP���'<"��~������j�Su��K���Lℍ�O�q�rH˴��B�N�A[��������.�u�v�L�/�����=fN��<;~!�e��X�c�meՏ��=�I��O�7����-��U�Yc��Q#Q
����3�l���vr8���<҇�׃��������/8�K���ܝ���	�B�|�_e���n<����(f�\��m��=�78��3���W�b��K�=5�$��t��F�E͚�O�[��l�dk
T�$�F���ϩ�ԇ@dG�R�?�+h�i骚��9,�|�]��y ��L5����`�g��쐟��c��G���U
^��ڌW>Z���w�:��	��"��5j٩=_���QZ8��E����+�t�cQ�4ꏽ�K��h���Ӕ��F@8�9+P���R�&�����H=8����=��L�	�Z��|�*�����ci��w�0�@ڿ�]i��c�2�AF�[u>F��EߙT@��n��uV��G���.���-g�Ll����B�9�?����VSH����8)}$	�=���Z����@˅�AG�˽�M
S�]!���̃��&�� �e�<|�v*�%S��SZ'���lT�B����k���d��&�Q<�3��×e��?���xty#�v��v҅~��PS2�Z/�Yt�t���`S�-<��R��� N����V�L�h���'�ءP�a@{KD }I�x3R��y�H�����fGet�h�������-o�FЈK���c�I�1��zU֐'�U͙)s������ EJ��,G�O��I�l���k%�TB{Q`���~�����Cl� ~V3$��q7��5�;s��N�vqz
�Г�^���+S$g�H�-MC|��me�A���[�a_F��W)�ąQ+��R�ObM�@㬈 LH��\^���C:5�?3�[�:���n�S��\~'��5��*�wY���
Av�Ȯ�R	���r�N^��+bۛ�$�O��xiJW&��kG�i�'Lj�Bx�2p����j#���v>6X޿C	�c�dp�w�2��"]W�r���¦����M�T������s�{��p�sٯ���g�B#�#Q[��NaR-�h��2o��1�!��(��X�>0.��P�{o�`��ș��+|#��4�k��kn�HP��?d�������&�^�ҷ��Il�-�����p�/_�@@ K�6C��F{�m�wh���y�j�}ߠ���qe#E�S���=e�?��7��e�sy��*;�K<���I������$��e��.i�u��H	�@����|R7�y҇�ew�̬@G��԰���[&mz!�S;��@�Y��:Q U8F�iVI��Ϡ`b����#�mЎ���*�_h�Z��&Do(�m9{��+^�n�������N��m�59����%5,8�xV�M+r��3��΀4�E��Z����/)Y��݄K|,������N/o *) r̉�)���]m�鈑"t�S]g�K��'� �za��n����ZK�	��3n.t!�V�q8@J��_�a!�6�dCr�%�l�
�i��=q{_S׷tw�]�S�0�wS�D�0g����}Bs
�L!��Z��wh}�К>���c`KI�f��6+������/�l %~.;!hv:r	9^�I���6�����(ڏ7��^��ܭHt�58�@P �<P�;xx�aIzV��p�,;Ql/����PV��۰��^_��?���
�/���;w���0��4Kյި��ʫB3=�����ygJinW~���1x�/��IC��B�	G���>FVYkN��N�1;#�ܘe�-'`�Pn�wu7�Ta��B�Q�X�?�
�����ũ��.�oT#�@�{aY�Ne7�-�$��6�4h��jmz=|h� 4[L6�cv��Lp�uLOhJY8�\�F��RI��Ұ	�׫<L��9�x�No��3��7�x�A8����p|1���o�}�2�⹮�]Φa�����"ġx� �x���A�P_B=Or��_���N�nG�r�u���g_:/���|qKN3�&q��QVm��]@ْ!�/��>��Ur�a��Ի0���?�B]���PU���+U18�K#{���]�RTI�����B���JZ�/���1j�������n��f�n�)*{>LފPb�o�`�i�<M�5��0����p?c�Ӏ�,(��\��u��i}X�w��V�B�%��bu/���N%��h�m.8�#Z�\�dO����^�P���S��Օ��� ��,�D���14?�s���v\���Җ)����Nf��{��?@�
.̢v۱"^�ȣ�:�A��vaw��S"Ĩ����lwK���LP��5]!��,-] {ki�cC�Â���{�k5����i��:O�ۀ�f���.�������7ܨ_s��K�ꄤ/GN_C]��E��J��.*! |��qy�(h�:���nmHu�d*|�l�s��	��{�!�����e���YYˍO���m-N�N𛽹�-�o=���+�,�����~ŕ �R
DP�)4ѣu��ۘ�!5k���#m��B��'>Gۯ�2D�dU�$ܖ���61����-��Ҕġ�	�^���y� :\A���6!��k3��4O*V���S,|��4�BD�k۽Wk`Є�W���4���H'���s�(W��)H�Sj�0,��~��J��w��������A�1�Æ�w��b�E��,r����﬚��b��v)��w:�iب�DF�,#��+v�c9�A��,��4m=j�������e$�F�{��>Ӈ1�5�I�%yZ�X�qkO��I�.�)HԈ����r�	��	[6���7�Ry�|��NYr��w�S ������va��C�M��'��d��|����؋(H*4)J�7�4A��S�vrkp���0>����Ǟ�C�F�c�`\͏�x�R�$��!�?�3ϜlVHǈ����?R�2dӐ[����#ݏ��̉������,[zU��Ių���s�*�]�2x�R�݂�N(��z�H��i���5Zغ;/�y �^1�L�3�iY�\_Wz�g1�R�!�L��K� 垻[��+*2�4`�z'��Gd5�T��Wd.2�C#N�Tr��2Ϫ���c��*B���E�=��,���b����i�[�c��B}�ߺ�ު�%��v^Yvu.� �gCü�����ʻ»�^��~�-n7%�N���X�PM@ݳ<��UH���@j�I�������"�H���e��.�_�i�ڌ���	��?���%n�B��-���k,\�O����2b���%��z��W��_/���? �;��� ����Ƃ��dV���h���z%����je@�&���4^�>Rd5�X-E9���K2'�v�E/2$�������ޞ;�֦���� �{��)�
�$�\���^��@�i��i�ߝۨ�c�W!@�=(&�:�yV{RR��A"g�R��/G	CH��gr\�2f��n;�	4T�4B��3�j�1������D
�q-,;y�j$˰z���]g/�8�B�X5@�r�6�n4�	�����Ax��P�(�iE��{~\��N�>ތ�ݏ!7��%�V� Y7�mY�ד��ޗ%��:폋��}�	^ǕA���2R�e�e~�4��V63ĳӐ��b�q�MRX�<Ŷ�����y�)�B�� {Y��.w����-Ws�#��q?��d��+p��f\����+N%<<�����.��s��������6CH�����b�jE݆������%
zz[ǈ�.Kp���:x[2m��t?�X%�����,Z�S�^�43������4�7��c�������N;��Q�Z�v77wH�S��w�	=r���ϣO!�jtxZՌ�9�I(pv�h%��
��]�P��>J��	,U� 7ϼ�F�/�L�G;,�O��ܔh����Bk��`�e����m�a��6�ɴ��l�����O{��v���B��L�z��9~y��"+.�b�G�I튦�E���&aD	�gH>�����a��ȼ��\E����}̓5j�,�Gu�Pb[`VT�(ί {�ߘ,G~lʝ�v]w)��MxZb(�8��Mm�d��v��9�� a�d�(Kh�=ɯ�5�V��ǅ����~��FPB�O��G�`�zJ�`K��y�#�����k|p}R[ZX�܂�X�����
��w!Ƕ�޽�j��b�$Z��:Fb��_y���N�W��9��ݤOoK�c��ђ��t���4�]�����|��|�:[�.�Bָ%�5v�`�����ٌ�Д@�XKQ�u.ar���<t�`@�)���NEt	�����@��5�>� K6���O��ͪ��,�T��:�|���a����Cì���#�\��GΜ�L�	S8�y�E��Y�'x�[� H��C�����>h*�xp����[^�����3H�$��Բ��9[:�p�I���� 6�P�,Y�y~���v��/�:d���Ƶ�(b�ɣ��Ut�f��d���|MZ��:��w:]ޖ,m�5���~^��;��=�9�П@籽_�l��YY�M�ӿL��%�z�uVǱ\6��G�1��ɇkL �۾x5�:ar���C��tl?�����ĐY����+���\{�«""��-{��*�d��x�j��߭�@�:\,�fnך�Y���V}ִ�mw
��O1f
�hC?F�:N<	�jy�x�-Ef��d#��@>���2w��1{���Դ��o�����"��O>��W(.��Fol>CbsEZ��������[����΄X[n������;��pA�nC	*��=cL���������Fi���:S�.Tg-�P�;�dɧ�/$�F��K��Ԝsl��t!�v��Z���㼟�Ψ/����M��$$C�Q�P�Yw2%3�V>�*����h�"+��@�� ���B����cU��v=�����(�9I0^z��i�b]�U����Mk�m�Uj�N��
����4��� ?�n]u�:����h�b���yd��m����`�}拌�4�Uf�_I���I˙0�	������_3���T	�N�W�w]3\=Z��J>
T��P,F�y��/��qw��#�E��ꚙ�� �+��t�]�gdݭnr����^��>j�|R�TasG�A���	�ay�g�d�� ��;8̗�B�e��~�,�#n1ߨ����m*f�! 6�]��(�ht$���yҗ���{������:>R���3��i��$1׋��ä�CL>�nV*�ٯ�s��@����$.�5ǥǣ�Z���9�$+�(�ƕ�Y
���0�:��#\��<i�ە���c�{���_��ҫ\j����P�	�o��ݽYJ��LDo?R���s���VV<:+m�Y��U`��������U��M16�k���!\?R�3�`�#Z�U�@v��;�ɠ�����Y��ŴZ&��$_4+�.�$̭B����E��Î���sCܥ��x�9��ÄXnA4N��8���.��~�=�s.�D�o�˝�u����I"�-����B+��}O.��c[^X��N4�̩j��*��h���A%Y�C����m�JLN����p\~Z�2۷V�Oc��B�jp��{���`�[8x�k�#��vI>w� ��`:Eb�3�����4��Rb�z	0����s��Y
��0�W�6݇�2uf��@8�rz��w+a:�n���^�����7�C!Ld#�g5&lj�P-%ۉ^�K���;�d�0_��WIޮ����bl�6`�y?h#��tŁ�(�a
���ԍ�o�8F�V�bLf�`׋_���2*�E�?�������|��K�.a��Lѷt-�Y7�VڜR��H�2�w�Ţ���VV[�VeӨ�]q ���!�tu���nU�wr�xq���{���7�>�"�+�'2M����JN;�@��Μ��稧� Đ�Rj�OMu`�x[E�@��U��!��pV��×��A7��^�h�aB��/��s�#��4�6s�6$�NCP%8��'������e����ʞQ���𾩑�u�	�UΗ��h����0L��;kH�=3��1+e@maYI��*7c��U���ď"�eC!�*%[��R��.'���+3_F!2'ԔՍu"T�� U(`��ʈ�-��3�8H3VV�d~�����Y)�����/�S���<�LU��Il�|�3{`�u�!����IY�I/��'+\<��7Ґ��U'���#C�F%�G�/�ה ���e
@?�+"�F�rψ�m9L�"�z+�&�n��V	�v�!>k�moN�����|��қ�������.�O6�E�2�U�3Y��U��R�w���?�{$�(����O���|�h�vO�'=�(��*�A�O��)��!�=��M�
\BC�������	��(�Jx(�os�������� o��Gc6煄�E�����cI��U�����=+k�^�O����R�<����v7@+Í0�8��g�͊D<p�A� �c��\�x�f�uL�]7bt�T�>b!�O<�q���3��=��h0��k���ɽ�r/H���=�t���@���� �Q瓳�J�����$�IKV�c^��_�_~��8�����[)V��M5VbZ�� ��f�)l�=�V4�޴�U:���'i�R镋ն�,0-�Hn"�y�5�C�$6D����D��������|����GU''7�۔�x�Yt�w���%NNౚ��02�pU:4l�Og�W��[���Ϩ�����	.�����̊J&�~�Ht��}�vC3�Ue��L���%�翽Wa;QըE� ���W@0��o1	*+cѨ��&�^�j�znU3�2?` �Q�J�n���`��1�5�j;poU�l_:��Y$������փ�j�B9�/<��j.�A:h1.[I��Z���&������B�&���EJ�T	!���ݲ#��^�bw/��RB��Q�x�Yj��A�j��e3�+�oH�;٠�������t�C��Z��sRK��l�������dH��3�t����{背}$� /�|%�[�hw��l��r]�|����ϽSC�b?A���F�)dqU����?�w�BE0�
g5�,2�<�*S�~���y)��D��<�d�,U[�v7
ڬjO��S�_�NŹV�@��6�#o����C�9/����x簶u�k�̣*�Ut鏽��-%D��N�p"ϩ�!�MNtEڤ��p'g߲͙���Yѕ���5Os�ʹZ�XŘH D,�Ϲ3e�$!S#��C�]���ؒ�>,��
�E����@ߧ��hX�4f=�@\�c�9�����%N���ѫv�+$*��a���s3��+�TtbA�6c��%g����	tg��T��Q�3���}n|4����q�+�Mf�5'�ę+���܂%�F�fx���!I�|j�HH�
<���Ӯ��OC9�J��K�T3VE�M����gS��'�s]�b����q0��&�2����ʯ�qy$��5'��ޘA��2�2��/ub����?�p3@x,/*��JS�gc��p����b:y\�.	�A���Х�\]9
��ĕ�cʥ���-�CO���]�T�#Y��;w��a��]x�0���er��0{M��[8�2�H|x�����WA��f�A,~���).(�4��I����>��$��!�]!J�{�u���ǆ�����v�--��T���]�u�v'��f�4�����Q�H��}���A!�h�!�{‏|ٖX�]_P-��~*�3>	!�*��NQN?]��FǶ��0a���
��������3�����j�Û�*�\�����;�����]lmN���は\Ҍ~
������;̆�N�W��=m��J=L����>�i(3�2����=��1y�'��R	e�!���U����evW���3��{˪:�!��ޢ�}�p��6ٸf�E]�4�c�>�[�R�^�;HoM�Z���Dg�1���X7jЍk��j]�.���Ʌ�e�g��9*s���	5��.g������"��n]��|U���"��1���H�tn���D;�����z]J������16�t��<��;Rx�Uf�/��3[�V!3��j�D�kl��ϗsO9J ��tY�?}�]��p4�+AT~
EauGmg?]�_�I6of�3�G�\�6;f�?���A�\�Np�`����ef�+$���T�+�`��B&�%}si�D�����="f�?K���
����
�yf>/�s�)� ;N�C�ݩ{����}|�&J������]�X,�>
"�M	7\1�n��kL�����C�0ͺ^�^�yW���6_Ci���V4�M���u0�N}�[�/���ʮ�0̧���/�����ݛ-}pSy Q��F�XR��H���NH�'�K�_Պ�w�a��[D���N�?w���Zţ�u �͂��� *z�@)��˦�6mY)�A4E9ј�r	�at��n��p���u�ݍ0�5Gv�'�\�Z����;5�mf�����Ҵ��L@n�*<������U#� �\� L-̂\9��m�u�+vemKu��׻Սq��`&��s�p���CRFV&����.@��!j@�C�4 c�=wk�֎���m4g�UTd�q�z�t�������M_v��k��q���R��F����G)P7���8U��9���*���\�)��ٓķ�]���gJ�ƌ����R#]?������tc�bzXqz��.޷@3���Hp�j�gw91�1�e��,WC�ܖ���~ƕ��O��7���,r�G�$8�Kp�kv��\>�?Uò���TR���uq:���M�lY�7H��'-�kj�ť��,�g.�o:���zw���DY��7�ڸo������+�:��&��������O!�3X- 
�	����/���(\�W�r�3�PCn�H�����5,�B��SFz�^�S္�C����'Zcʜ�b�IX���^N�	��Ņ[((�a�3��͞�X:���M�eq������x
(Ab�ݹ����\D�/6;��x�����!B"q��.���-��|�m�	�����p�=k뷿6�.5ۏ�Š�����E��v��H��Y#{��vX*30��1�d��|�p�,5J���9�K�l�7i]��(�Z����BtCм����.�Q�~�tc��f/�".��d���&���{�&��cSnzCM>�S����pID���R0���wߊ��U�Ǝ逤d���Z�H���"S.4I�M!�� X0y9l�2�-E�������˛�J|�������`�l�=Q��-o c�~�e�]lc�]��7Npf��f����. ��^ �O�1ֲP�Q�f�"q�����PZ�E�	J(M$���a���?{EO[_�s"c:�����A'o�n7�&9�8��!�P9��?G��pNy�>V`����K�F,��e^a� ^�UN��#��}�c"����z�w�/��W�Z9[���@"|��.Qƃ��QN3��Z���m��❂����Aګ��s�����l)�J��qd|d$�x&�5"z��D�ۓ�4��e�\~�{��Tֳ�;|�K�k��0��ӌ��-�P�$�����7�Lgj)���j��O%k�^�[��7��ko��OQ~z�@����^TLk�֯�@�$&(9�ɬ�*�f`�\��h�&vo+�Ҟj�A/�Q�XKk)�Kg��A��B3r!��2��w+BeR�s��2�*�s��-�V�[sx��z8� �}"�sQT����� _1>��@`!05�q%��3�E ��m���.�3!:6z�`:{=3�Q� ���L������1�q7��GT��/�b��7�f����|�5ʼA]���͈�/��qt#	��ZgkCH�4;��Z��.:����)�g��ͫ
2Ib%���i�U��?�):�rD��"��؀)�M�bp%��'��h�$��hY�B[-���m��$�)�<Z֦͋� �B}���	���)]��,�Ui��W�{�x	������\0�m!=w2��Tx�)Om���z��^�2�ջ�lm
�GE��Ў�����a��%�I#�5�YO�8\�.���~�_��2�/�bm�W�[�˰��i�˪����lrY�
A�f���'���T��u�LH
��K3fu��z��5'�sqگg��b� |���R�Q��>�Z�j��p�>ڕ�S!s�����9R��� y��n�]��D����H����X���e~/$ƺ��(���3�Ny] �����!]G7#!�K�Lz�
Id�D�����}HA2I�"1E�-�7E<+��Xx��])�����Fmŝvxn/���ɀÒP��OU�,1Z�F1T����zw��[��[	�]q������;f�3��k��f�������G�S�y6��C./�3��tW�k����|ŏ
�5�Y�3����Q��N������W�k�[,�f��J����t��ݔy��O����.�~�"_n�5G,��o�ٝ''Ŕ��տ9�BapA�C�|��J!Rnv2 |{L�+�P;�GyP�8N;����锒�HL�N�o)��t,�@[}��(G��Q״�A@�2f�@�Fd����U�~�(�����RW�)M���)��+�;�G�>n�����1��F��N,�e��nX�-p��[Y��{z�[�U�����s��f� ��F�2L���s��i��,���虾+,;��t��c]9�`Ҝ%��YɄ�����o�;��	("�U	{����H'�$�3�Rl���(ĸ=�5R��WO��Pτ��Z�����}�i`�1��혌���yşFM�
6_R� ��B�滈����G��ԑt�nG>��z>75#���>�Ͷ��V��3�,�(�������i45�q?� �c�xWV�	w)|Y�VA�f�R}���D��i�SG��2ε��$�I����۞9�_~��(a�Eߜx�g�����1����↜>C�? 3M�<>+W6�p]���
?/�ۋ���^.��Cz鮎4���m
�������gz�(nj�!�0�D! A����i/ۜ0Yy_��Y��? �o�.@�й���:��t�l沕F9�
{_�זԌ�>�����yQhd�+�ۓV"'ͯ� �5�9a���6.y����a6sÁ�9&M�p�yAW�m!�?�Y|��	x�Ƣq���������2����}?W/-/�����R��i<D��G��@�C�Fc]�q��9<M9Ŷ#Ҧf�,��N:��jt�ȂT�i[w��������3'��DBn�L&�#V}��b�.���4�N������/)��� ,l�]�GH[?��(LOѺv��,���bT��� ޺���!���s��ʼ��d,VDöt*r�o���e>��ǫBq����U"2Y��%���':e�RL�-��[��Ǉ�q�D�п�_�����^�L��J�k�ȠJf�'L�f������?���5:��|�ʑ�Yx����*�4��!YV"�|�<^et���"�"�w��b,��-lXq'�����7��&���D@����+T��5�W)6�*�36��Lg ���eOQ��X�H��F��{k/�h
�f�wo�ca&���.nӮ1)�x$��wEi�`�7��1$� �H7Θ��l�`|�^�p�
�bο������û\_ᮚ�s7�b^�x�-�y�;.���{�l�ȕ���c9��J`��:N�a?������?�t��y����ӣB��'��!t�ug�F�з��BÕ��K^�Z+���GݯG���+��I�؞<]�8�� ���:���3;s�_c~�7Y�2��Iw��|��o}�^�{�u�+�-�\���b~\	d$r��*����j�=�Q��r!���9.t���t��*reK+b[��,^�,,��Z�
wT�d�Vεr����g�2�nj�_,Ur��*���2 )U��fR�0O��'��u၂���e&uy��J{e!	���d��m4��`D�x���=�և��D,N�:fE��oܨ��l�b������V4X�dY_��l��	��[P�{޲�2��|�A���c����;�B�-�қ��Y�T|&��Ie�������n c�r%�SR<�҅��F5p1&$��/�� n��~�����(�V�C�g��f��E����X��7U���N�49zF �ל�;n����Ќ��칻�UݸZ*q2����^.ޤ;�䉤���g烷
�5%�}��Z�=2T�
\R���s���
�ބ�ܷ��$(�G���Y(���.ks=Lk�`DϷY:'Y�~!����~�b�kS��s��B8���na�D!��W��+�`�ϯ�z0)�ڐ��c5ʘ�]�B^�_m���u�Y6C,�P9�T�S��ҳ:U֣㍘ʡ]�`G�5��:�v��_�e���d�6�N��c�é��#_��5=z��㻴�F�]�Y�0'�r14�|�&s>�l�]��vr�9}hT@90�ߧ" ���$��^~�c����g)�r�Nժ4�.��iR'�(P�������7�@���$�#��Z�r��H 3�oFK���2E���.b�Dw��\b�~�r��=�����d�4�
��^m��G	RQ���k��V��]e^L�?�f.�=�v	s��w*R�邆*v��M��$o��:WwKI��j��]���a�nu�ɑ�Y��jj��8�	߅�Ȧ%�r�F�^I�z�R�Bf�V�7��N5��V���+���+oAF��`���}��٧�{䜐�{��C"���?f�=;g=c����u�8�K�*�(����v3�W���ȥY_�C,�+����h(�+'�Uv=��N3�~0-�t���f���|�i�ZW�7��c[�D�l1ioC����/O�,4�S&�z~��á0��E*y^�{�Bg|��W���o G���e���m��ǐ�|�)r8�]��0K��	%�n�������E[^'��o.��$٣܏`���hH�!''�r�7f�,zakJ��TC]�R��e�=<�8��.8���_/��'a`>T�Ƨ;����TL�_Yu� ,��b@\σuc+��1�������eGeW��M�|�M�>��u{>s���U�b���w���?��:o�/�xX���W���ߌ+���7��`�y�JH��N@"�jt�2+�*��Ӗ����]p�hLzJ5Uԑ_Q���X����C-�L�FeB/���?��&=l/�(��Lgyy��yTd�����/!�pP��w8�Y�&D�j��B�6�pPN�cY�������~�ԇ|(FS!��L�`9��z��2��z�}��q�7?��K}󰏋��x�m�0�����t�9>��i"�#�� ����Q���m�T��a����^c�4��#c&t�SK����A��=zc~���!/��lbb^�I��C����f�[{ͼКҔ���UA}��>�q[(���$��pY�@=��Ɯ�oF����R!P��a;�p�C)wr�`+F��^���f�]?mhy6�Th�!v����-9�Ea�R�$&�����^�vX�pH��c���-��|Vr�?�"y0>/�=�06�|��F�H)S�D�6�Ơ�2��*z�)K{�lN�G��G��}Q��*+�e��y
x3̩I�.�[[�o��&����P~���?g���@��9�AR�3�aN�G������ދW��K��NŞ~����$���z����Hܿ�'�N;KV*Bno��?�:����:g�-z��_�P��	���l`�Z��K5�.uT�;�u%Z��u����M���b@���g��rZiZ���"v���Y��������!K<��������U(JU�����$��]�.�uZ���$%v΍�r�*W��Φ���^Y��	&���Vf�F ��܎|�	و��B%W-fl��L]��hd�@�7d*a�Yb*8X��=H��$�ӊu����i뵯 �^3:'31�t�)3�Ҥ7���U(<����D�Z��ۨ��5�p�'�(�̱�Wy�4
��1�0+k��n�f�F�+p˪N�۵��q�APd�tN���H{5��V��ѼMdE�n5��J��jL��m��Ӓ
�{��Y�Ͻ*�*�Mb@u��k���1�����7�=�������ㄚ�M\��'/�^�׸�\��ض���MM�
��]u
ai�pO@���8Z���j�dQ�x{i���r5�n�	���6,�H����Ԝ�2�}����v�h�f������Ė� ~�v)W/�$oQk9��	;r~��x&0�8L<MK��Y,,U�U��Ѵ�� ��r�,��H�@*���.����1�.�^�1.d��j5G�c^kZĢ��g��is�+��~�T])�\W^�"�.���=���Ek�j�!������<��VM��Y<�]�6�#��K�$hg�� ������o�FD`N.���R�H��ݠ���'��g��zG��j���s=�]{����r>���g�)��i�1y�� ��F��VkS5R��k�e�ju�	�H�H�>#\G�=�Ǿۏ���J�_�Z��: �Ķ��/��D)�w#�sp�v4���J�� �s5r�:˱���|�h����
):�j�+�)[<_TR��pA,����;���0e��(o�$� ����u�����/���t'\��G7z�Z� �W�V�m $)����gܥ@ı<�>��{�Е����*�ʗ���v�\�i�$��d�&̂�z������L� 4��m���N�e��nü��[PE?�c��s�΂��؜�}�����"�Q���2!a�%O;�p��[�1t��`��At2.	�ʂ������2�`/~+�'E�T��?K�=��i��=" ���� ���%�͝9ta�w�3{~k�D��F9"��~�x3��d����m���[5oM��}ܧP+�rI��xP4د�q@�	F������.�6)��E����!^ `e7C������0`@�I�r�q�<�M��P'6�~���'�!�C�I���9���S�"S��R4�I�˄B�ӑK0���9��� �10����i��6��s�O� �|��.�.M��)�g�e*��l1���F+{]ԃ�aИ���[\��={��Q����r�T�W�9�̐����#�S�� ��,T�\�eyn���I*V����7�dvX�"P���I�gO�"�}#:�e���<��9�W\0h��pMh`&2���de�~o+U!Ҩ.��(�Xc��":�¸�Lh�D,n^O�ʲn
�m�x��h���d;gK��(\�(��f\�c�K���$ �@gĪ�_x��+k"Ql�����*�"�E�W���z�<���`�=w�5��r<J�\���D?�I8�\���zPr/qDY����W+i�au?u���JG�oB�N[��#:R�-:�����R/Q x�̗�-|�ͤ����7E �J�E�ދ�t�u� �������]o�W�t����� ,1�J[h.d+� �����GNd��NX��ע<�n����F���&:��fA9=ҵ[�f��;���g���\��NX�Y�ie>��L�s~��VF2��Cg~�/U1 �!7��پ*]A!KZ&�nk��A�gC�1�2҇��a�|�\��a�x���V>�u7\/��8�r=q���ܞc(���q>g ^�O�U�|u�z�$�Z+�0�S��C��L�9�-Ӂ纺���r�o��h|��tHD3��!���������ij|AB��+D��8 ,x�����|���z1	;1J����ΖبF��$�Bc��ua�����;�,]H��8\v�
*2���n�J�7�����]��B�#`��ڟ�I�����żL���E�Q�1�������_�8G�PGѓ�:N@E�>�_�<i��r.�К��o��g��&���p
D�Pl`>ݥ�w��ޫ?ȥ,���i���=_��%�G��J�Y�So��ǖc�ĵ搷>�Σ�f��\EE̐Ƚ���3��(���{�Z���/��J}{���:m]��ü��A�>� S A��bk�W�w�J�M���
G<xӮ�sNUĂB���8�A0���^7�R�ɯ+&�_~�9��YmW�@�����ȥ0-���a�N�~F��Y�5gw���_G�@:w��;��������	��% G?�j�+#�9@ �>����c(܄�KpXF�ˢ^�>���|C��e$%8T/z'�.��x!��!�ӓ�-q}'���98#d�=N}�ZR��6m�&ث!��5j�D|�)�h��!�t��wNS����/�Eպ_W@M��l������	����g�24[���[��6d^�F�/\?����Y���ځ3F&߫�=�!���`'��(�r5��=�k�<�c�w�S%�#�4�c�uG`|��sv��<˫c���6�t��Ō����� :�'��	q����iq�6Ѽ���k�3�/�V�YJƪq��O��Q�d�Ϊ\QvoR���=I�R��X�I�by x\}[W ���_Z;�JNgdzL֞	7gb@�`���5��W�i&�}�=u)�����+����d�-�63���i�}����g�hS0{q����e�a �um++K��Y7�T�oua:&�����b�,���T7Ԯ!����y^FR��h�NY��@Wr�;ʻM���|(��M��!�Ey~��*�}<�ه��{�0�B�@�M��\%�,���^H�+�(D�C���UN�6�;�'fNS�(鹦��}�?�w$���[1����u�d��]��H���V��*��=��T!Ez��T��MA�*r
���x(E>���K��'�z^Xj5
���h�v�K���|���>N�ʼ���C �M�e�nk��i`�C�sjB�A͠�F�mݝ��F��d!�O���O7t�LP��8����8rT�f#�x#���n?7��L���^Μ,�}>��*�C��;l��8����fF->���o�f�S���Ţt�̼�Y`�^x�p|im�����4��+�@ƥWn������4�o��01R�B��K��Xy���"MiԘ7l��
(��7����T�12����`v�_r�WynQ�J���a�G�=��W��
#�p�$0xϏĬ�������i�a�B+�@���܃�#�~�x���^�
/p��w"��kT3� �x=���I@M�l��o V�c��GjS����{D^�\LcI�4.wK����,��{���(H�E�V�H&�:\2�n�809��Ex���ڈ��/����7��b/�$i��^i�#�?Э�l�T"��J,� ͇wU�=ۘ������񺾲\袰��Ro�Ֆ���u}�.54N�v��4a��9Iwyn����a�h{й�F���W���Nx?��+�(w�/|)�2Csw���6�ۇ��p�?�����&F��nI������:�F�u����b]��Ds��$Ti���J�-z�'H���y�⸎��^���{7X�]q0<۳�>H�ܮiW���P��P8�A�&��H6�	b�?��1pM0D��/�x�*�):�(!�\��%q��<��Y~�	d�UeL3��Bك������!���δ�'$��ޠ!_#�|)��{[�S�G���|���X�|LA�O�e�j�ӄ�5����癑U��|ގ=�h�T�(����l-g�0⋨�Pm�w�ݦ�cԱ��ߒ5O
�!	F*��¤��O��Mr��U��>�<�`��Q�)������H��=��9����&N�����eJ� ��`��8TE@�����f :�h	���ʹ����q7�U��o���U�f�9��-ZW?̎� �������RƜԟHM]� =Fx��e�V7O�Ps��YM&Y?��N�ޝ�m�����V���B9�)��R ���5Gg|Gcj�HE#����%���sEǿy�V�~�#J�E#}���RR୒�礥����2��$�X�@J�2�8B���}������P.25E�}��JC�����
�[�R�~�\��XŬ��M	��W��j��2�g�%�}G����<xbUi�l��qJ��D�X�R)�	��z�hk��ߎ��sBО��Z=oby�k	L�i��H=y�H���ڪ��r�����<V��U$�v�w���H�����sYYB����JT�/}�ݯJ4OQK�yݪ�$�@ |�$��!�h���\N-r�Z7��˥U=��eBh����=3�3,#�-]oz�1�!1�4���'2��Ţ>O/��꣜����BI�Rm!��|��ӽ���^�jx����&�QuR��V��RB�^O�J���؎��c��>��	���ˬ&, �Fc��DCMDI����/��띝�?�
3�by�4#��'����B�_�JyOn�P��O=[ �)�s^o�x���������J�M��M��.�+nͪ��l�U�lC=#܇��I@�)�1s7�B����3�Y�ܴ�
p���؀֮Fxe׍�-��c��D�� X��hm���`�Tn��ą3�>G�J�/i�P�q7aK�6����ϑ^͔�O�Hw�u:1�v��ܦc�+���Z�O���h��Bk9�JEG�O��8��P\���!���(h�b$��Ku�6L��%f����˝36��t�TQL�=�>A9��KlD~��C����sy��hpH(�,���r�i��,z���,�{�[;�Ӛ�Q{�%A�S[	�o������\�n	�F�`���Y�������*5�8��p��9ٴ�� %�̾� �"8��]��?m�@.��
n���V���T��T,"SC�5v*��E�.�z]H2�+R�Ts�;wt}ė��ޙwC]RR]��57ha�B����^�޸��š��Z�������um��N���k��#U[�����j7��̺��xV��X�D��_�\<믜D��zK�M�r�\���ڭP35���W�-��?*V�ٷ�_3��5r�h�,����訅��"(�昋N�K��������M*V��j���t��2��
�&�����*��l�u�yu=tG3��8:�vR_����R��?ʼ�O'�F�S��a���2�4R�?g�#��M�,I��S	X�o��h�%�K�֜IN����ҕ-�>pa��@�+$Ж�H�[��d�����,*ˬ� \W�C��w#�$iyC (�<Ih���@ٸ}O�b������������(�z�y�S�8�AC���%CQ����7A',e#�h��x��}<l��h`��o��Jձ}�~F�d�L���۴.L��fʫ�����Ue��S�+?~ ����qI�?�~8�
 ���$��'�s�8�fs����������|��]�v��	�e�}R����d�Z曾
���m�ej��7'C�e�'d��s�3� 꽒@pba�Ҋzf��_3��,x�$��ޫ)��^u��r�@��xI����=�mM�q�����XP�C��Dt��Ԑ/�c�J'�W�4�ʋ��k�� ZA~�����"'�)�|�R��{��$����|��s�޵��
�WIo3�W��4hA,T0dv<E���3C��b�+tU����-�s�|ל�%����يɜKY�����).ߙ^�BǺ>�l�g���R��6ߗ�,(��G� z?�-�8�Y�*ZOwa��W*�1���S2%�{_�m7k���E�!)o"����PZˬ�ӓ	�J�b@�U�
��6�;��r">�n���[��UyTfQ�X��9@�A`��CJ��Myyl���ͳ�(�u��*a���݋�՜�����ӣ|�� Ր���w����򖰆3��1����r^������M�,�Ő��a��,�~X��+�NH�y��1|^��]�Ri5X�����uɯ�2���X��^l�[�`-��J���	��c��E�h�ML���#:�i�G�����,)��颐ë�D5a^��D�T��y�.�j����ij���K�����z��ex��7aJ�4H�(Bi)|��M�b<[�%�7`����>	W����t����I�?\~yBޜ�>�]Gm�d��S,��r�� 4-�iQ�S�ͳK�85V!/�����ؚ�1�KB��>��$���]?\�sN�X₈i)���J��9
�i��RX�
�HJP�$ܜ2�j����u�g�7&C@��YQ֗���W<'��ߝ|�(r]� ?³�/��Nsl�靝 ����>	5�p絙�a!�W���9-c}H�����e��F�?�޾F>��C��6~��`�jw����hS7�p������G���[���-�k�iL�k",o��ǓG�(�F�qB��@%h��l`$��@=�s�e9H�z��B�1{`�B�ᤝP���=��d<�1���h�˶2�6���<i�ɀ��MG�d�`�O�3�龶��o�ֆ�!J�a��i��A��O��Ss:2�(+�I�377 !�����m�,S��^�����uv~��R<�`�^7�ි��s����3ە'�k�zA�n�m���a���� G�g�eC�����H��N2�	�;�H�����>'҅�d�Q@�)΅�f��G�F�̤�27'�Q��쏫�9@��Il�!�����j~�Al?��(��o�ݐ�pG�Zz�LA���m)�81�<��1��b��t��,��[;w���GH��\�'��6�ORoB����6���1mxR���c�E�[_S$�0xH#��$��Rs���\_�^?��j{�Q���G�6���A�#%� Z�3�`ٺh|�
�$����z��}M�/��nwf���ɖ}� FH�3�(I��o ����c'��;���'g�7&�V!Y\�/!��4:���x�0�!i�nzN�-�x�%:��D ��!5�Ri^?�OˈY���8*���0�}?֛.�� ���#����L%$�}'K�o#���ȓ,�Ch_
��ss3'��Ԧ���X~esc���"��w�V�7�i���a��7(V��R�	L�W��
& �-���3��?P��^���_��d�w�7�� gt6^,~�D���ԁ�� q���4o[c��dg�Z�T��2nd\��7"*��<<�L��s��y��a��Z�gZ�&��s��w�j%�6��\8S(Sk������}�df������Bу�!@��I8��g4,<�d�	*���<Q�C�^2G�Za�X��'�,�2����_�|ڌ�qgk2r�ܼK�/��U��0�V�-,aUo����(c�nQb�ox�������%K��0S1����: U�m��vTt�F�V�7��ַ�������MN���<	:�1�)�k���p`S1����l6O��0��u�"��K7��8���q����Г���V#$��6N�%����4�.�[<�rީ��V�7`��\�J~�����$ ����.�pR'��^֪����k�:;H)k��9ӵ�,Q�T�9���{wC<�#�I�7�
�_����7p��Y��W���%MQy��-���g��� ^3"�l�x�B΀V#��C'^�n�l�7D�rH��y o�g��[�@ôEȸ�� u�-�s��!�S��d�*CqK�4ηqR�|��@��tz�M����U@SE\�ov��k�f�;�����wzJ�u�+|K12a�u�Ux&(Ʊ1����O���і��Y����IC��ௐ�S෽�ߵ��B��!��t�R��<_1N�>Q�Q�� =Ǫ�U�=�ŰR��E�.�M~�"پ8��$>��[������b���~4RC
�:\�,���9[�1e}^���r�0�`�7 [��t폙��3s�
V�P��d*�Ȳ�{<��|�%>d��3'M���T���oA6�K�{e���Z0�鲬���5�����C����E����A�����
���XG�����N�����j�����\Hl���ׂ�G"	ꉿW/5ώ�C��U�{u�$paʟ��o
������.¡�~�kyz�c9�A�\���87}3�1��;�#r�ΰ"��:���:Ot0���7��V����{'|�>O���8 >��{uf��]��q3\J��lXF��Mĸ�����4C/��!�gA�����σ�5xU�k�0�]�3�_@!P�n�� �-	V��K�f��:�%�t��K҂�������r�q^��U����F�jj�h��1(y`9�8Ui�D<��϶o�?�s	k���7u9�Xn`��í�hP�f�b����󽨌T`+��9s�r�$�K�����p��X��,�sj��O���1��r�đtVW��>�8��������S��_�G�R�������K������}����|���l���V��7e��o�`|P'�f�s\3�0���"��hU�LtÀn��/q�98���\"Bt�E����p�����h9C�_3\��i����*9t�͠I}_D3M=k[_�f5o��
*hB3<��*L)tps)B�O6:2ޛ�N�7w&i��̗L8�`}i����T����>�n�8 ��:��%c;�n��KX�6mn
dN�~��%�(���@_L�<Q��|�_���?�Y�-Å����w
 >��S�|w��x�"6���0�
}�Q}�RlyŒ���V�r��>���2��廇��p���G�)�[X�U	�����t#������G�7�#�ᐟ��gB�.O��u{E;�IAo��y�.��r�7�$�������Q���>fuk.��zr$�
a�q8�Pc�z�7��ɎC���ޑ��(����tjX��sq�m%�k}0��X����Fe/��8n��Kf�m@�ּD"*�Lq_�?��=�3L~J�@��=������C�=�<s�&���.;�#f���Z8�^�)ɾ�N�ڢ���/�����:�0�?�-9KJU('q��?$Qo3��;5��,�4%m��{�l����ܰy8V�Z��NӃ��xX	b��L��[�»{S(V2nӟGb<��R���aw'ʤ������H��<�[%�u��O(���_�����MB��R3p�����37��'
76|���C���R*��T��׆��� :�w�;/A��('�2�C���M��s�E׸�`����;��kV���?�	�4Y�S��S>�B�Bl��gny�+(�[N)��а��v���mc`���*�����Wۛ��\L~��_ꇔ��f`\:��kmdx��4�OJ�׸~��� tD����l�ń�"(��{���B�H���R�oki؜q@���. �w�;�*0���E��R�:�zuK1.͈�g�猯m�i�0qs�6w�M�K+w�ߑ�>0es?� )�6$4� n7�i2�((�	��r�/lfvwC�����O�]����D�tH���(�x�yq��f_ b�&�6���hf��|pU�q�w�����ޗ�ȝ�i�XF9���U2�z����M�O���M�"����F��O��s�#�M,=�(��ٯe�/k1r�z�ou�i��!7E@S�}
�_�蓻�Yp�fܽ��~����u��x����m�`�]���߼�i��7�ƥ�����]Y0�e�H��g��PX��Ǒ.S"Lvd�Ӻ7.�vI��ߍBM/A�0� ����>!҈��k�������e{�k��6$2����Z�o@y�G巟�t�����'�`�[�=��Q����|�<w	�K�9Ģ>� BIX�	H�x��tfQ�ǥ��Q�c$P"�ZZ�`��G�}l�׃��VD����\nL"��GQ~D/���"3�ͤA_�¬{b�l�L�?�y,�\O�["ۈ��|�GG�FR^�_�D�o�������'T�䔨�>�7�����5�%͖dƾ�m�ȷ|���v22��.���U��y�/�L�������S)]����t�+�{���%��,4���K\��H���̲{Hԩ���Y�f�3��A���J�-�'�=/3�"m+�2�+T�zu4�a�59��J>�W�E�Ҷ�ACM�rYY����9!egi%,�v��G�$������
�a$Z�Ig�@*��e��0,A���"@~p�]�LRy�,H�#5����񸰏K)5\���2�ܤb���@�-���.'�ݥqk��}�Bom4���G���v�+U�{�H�~$ݽ"��{[�,:'#a�PCE�z���[ٗ�Z�ƺ52��ZV����M%���!�OH����q���%C).Q��p�p	�>ߑ���	w�%K)�1I^]d�qk2��"�� ����-B�14tO�w�ZZ"���Ј�L���� �P>�{���n@<Vs-��fy+�*!�|���x>4�iX�b�?�؛㔺��0���55���6ڙ�������y(3F���3�mU������-R�_R6���S#F@mQu�~N-3���N�˓���4&����sS!�|T�^9��ض��h�"cF���V8I��ZV��6b �V�ET���ݯ�|7���~��W��B���A餲Z�N��g8�Hg�a�����lY]u-9ͺ���k��~�X��u�jL%�
G�?w��h|N���x�z$:v������y���c��N�i5�o���#�8�t`��������x�_J�j�{�|���`����#Y>׿D�{�>U�1�G��x�+aƾd�7���Mu�Aօs�����C��*�~��Z^A�#���f�Ś�Ȃ:a�a��o���z>���Ah�K�k��
"v�����ۂ	��(l���,=�ᆕe����_���;�Sf^�f���~��;�x���f�7������N����=4(�Wr��.YG	CR�:@�R%��]{�*�s CbH���g�_ۡЯ����#3��m^)'[?j4S��υr�gS7�5��P@�Ik^y^Tq+{{֢�V�9��K^���u,oEHj�;��8�>�x�,cf�%
5#���%��ueŌ��F���ƿE�v��]�	�w�)0�F����:�}l��Q��S/w�!�	�@ux�Z?����Ye#�7��@Ç�r�-2�`-S��K�S��!%���kɋ��6��o�軽M��#��D�������D�Ǟ��b$��Ԓ{��ޟ��_�@[]>���~�۴���ޜ�K~��']��r���K�J��4�m3n�}����R��<��a}�J��帯�5E�nMx��u���0g{�[% ��?q(^�2�x��V�)<ʌ�a������ƀ$g2�8�%���H���J� �!]�tB��i
���:`{�?	�����ӗ�zN�y�5��R��oMk�\�#_�N3K�{�Oh(��c ׿4�D��f�(P�M!�a��[��q�3�Zl-8~����s��Q��cٛ�$+c��.+�/�!F	|D�����N}�x�Z�.��(�W�?���AB��|z�x��iŎ]���vD� ��@��	ߴ(�G���b�K�O볩�lQm@�.��&j�p[D�H17m�%i��<�ؓ���|���.�>D[\�TsY p�����`q�2f����!;�gY">3O#�R_�w6%�;�]~�����y<9P���g�g�V��u�k���QQ#U3�����Z}
	��[f�B����H̅�&�H���+nj�#�1�%z��Z�D�u�wi��IQ�1ƈ���֣���q^@T��J̙s�gb�0���	�
v�)5ٲ��k�1���5��Jp}���c��~G��6��;L4N{��&�Ȝ�\H#��s���.�k�I��,�AH�������7�0E2�d\���[8H	oj��0$E#CU-aZ5�*��a��{�C�s�Y��j��0s/�{f����`v�\-Ϊ�\��֚�K��/���m�SҒ���<}]�JtB��z�����z��'o��i24�n��$�D��n�y��D�و��k�fD����	�x}h��ݠh����>�? =��O����8[@�������9���8	�]pcG�0���.��w����?��K}/�8Fn�^���2elu �W��AN�����-���V�-qײ��*G�Te�=���K�o�{�:�zX~aQ���9��&���rU@÷�Ս=�L��fVh`�#T�F��p����r����K*�����P��4��q��}��$R��+ew:h=ǀ�=���CG��i�E���z@�5>�UD[�+��͇���;�SH�ڇKTa���	 �	Otg8�`�c�`���`���	Q���Jl�O����`�����M[a53T������^}���,����ȱd�1ʊ.��1���3N�Jނ���0}�r�к{ (Ub�a
6z��D��(A��*Z���:g��JO?[[��El7U�s/p��w�m�**+��:�f��t� ������j'��"�eGatG�'�����Ӵ|y��������F'H�|oAxJ����m엓�y��AqU�@���I��2�H���l���	�q�q���Q�s{�Mu�{��4�"�J�
q�x�[��%k�[\�<]A�C�	�����
7�T��ODϤ^��f��A�~��$�%��/���t	3s�S�I��".�o�����V���Y�����\��j��2�J��=`ʠҷ�Kx���"1>�YhVX^����by�m]�|�������'d���݌��/ȼ�K�]��l3܋0��V�Aц����]�~A ��1+�-� TvN���]���u]���L�S����]��p̥	������Ԑ79��M�%��7[�<XG_U��M��N�"1���6�o��P{�􁩷�b�JҬ&}h��H��ҫ�83eD���Wk<�R)�0������&�pR��p
2�|���+���膠�j�E��SŒ6�M=iJ<캈�
5XC]J B91	�kb%e�v�T5g�}Oi�]�s��~A��G�0!+7��,^`J)��Iُ4׮�7��m�6R'S,}�{��G�k�	�Y�
�v��`�Q,NW�TP���y���9��p���յbQ�#I'*���X75$a�A:j�N�����]*���j|Ǆ|8���J����7,v�b�r�$��@�f�8�Q��6u���3w
�ٔ��1C��r|jt���t3�g��#q���7���#�fn��"�[��h����W���v\JQJf���spO��+nPm�!Cr�%bFgOD�I�NL�U��G
�NDz@�j�sl����V)���ܡrM�ͥJvǸPRj���pxh=��
p�S�ɯ)�9�V�N�Ki1b߷��I��*��w�<x5Fo������SMŻP� ��z��D@�GS6	q��=P[�oI��,��b-�\\RY�ف�2Yj�ŨA�����F���c�(���DG���AQ���Ā��eU�z�`@�,ؓ^(22M���%&��s�L_=A�|�E/����K�Lw�|ŝ|�/�9��;'�����h�_���u����_a� }
8 ��~�n�%k�W�:}{h\���1�¢<}��
|�RT��NP�uV���@@�������{̄�
`�7���m��fmI?-F�9��r���K�>�"(	u��Dp�<9#%�^  �����C��(������}=Cdj7�9ӎ��'�s*E��v���٦���k�j��0~� c	�2�4l7H-/)�S���z��U���`|�r�Vx��q����%��Đ�n�pK�2�D�o$����U�)�s"3q����6��a;;��ՠ��n悝�|��	�m6������Zp:�����/b+���ݾ[�Wq4�!��74�3��t�c��酚X��Q�l�z�o���h�5a�JC$�Q1�����I�$/��WW;h�}�c,��-YӦ���I� 2h����PV�c��˲9��jDL�U�߲v�HD����(�.k�E�^^x=�~\�8�:�u�È������"�Y�D��-�H#Ŋ|�=��)�^��*������sf>�����:(;��,𽸔붵�G��΋\Op|S6"}�&i�N���aBN�����3ź������C��&�V���&��L��K�!��`���vWx��r����vT��:ه+��'��5�C�E4�b凫o�A�}���1_�(X��bMG���p._��J����?���F&0�UAI>�G��{�w��#@<)�ߏ�Z��E�f�JR�o�A9f�6?�Ofz*ڕ�Dԇ�}o�����|��#�KQ��(1vy|����]���Z���2�QM	�)�bR��ԉ�pX:�2z����JƧ�<`�e��~�@Z�@=���7A�
���/S;�M� Mab�}�h�#5r�@j���,B�U������e�ч�Hb�����J>���[���#��p��%����B ���%%�1�88emh�n���B�,?�t~�p&ݞR�J�����v% ב)����5���'�/D���������]�$4�[�Sg�gq��)��\���[־!��WѺ"��lJ��1��!�U+�!ZtZ���C:�%�\�,\��	�"	�#�-�5�w#%��/D�g�V5���{�::��%z�����8CGr%O��H�kN��_#�E���X��Vζ	D&�6F����zL���~��|A��,Y���b�qJt��ƛس?��:�t�}�?������Ì��k����O9@���M�h��y&��v��O��'ڜ8 [X/�Z_h"Ε�xu�ľL�!�������UuOm�N�B�������N8%��'2Ͷ��WT=,��SM�-®kH@(I���T�t�a/��ؓ���~�W߻rB�+��b�%��I�u��7n��9��7:�t�Rzȓ�.*�s~��բhy8��<��#~HW��] ꊪ3*���|"|�Qn�=�(ʵ�Tx��	��x`U��OP�l|~���>9E�O��#V����������D�eN�B����A�[DK�%g�/pa�/Z��&H�iH��YS��~Q!1�qs��ː�A�?ً��%�@�<��=�ɼ��[���׺�v3C����. ����h�����Eت�F䋃�O�@�-��wN.�EippZ�dX#pR��x��a��D�E6tE�3�U�t��2�L�ּ�o=i��8� �B�hX}@�8����Q�+'\�=5��&�-���)jw%n���[e��o�0/uϢ[4ϗ+%:Sܐ��Lax�h5Z(�݂4$���ݭ�	q7��L�G��0�?�vn��&|�~�9���� �G��R�����$q�:�Znp �[P�ŧx��᠏��/���i�����%���$�%��fQ�?�����j	�u�E��p��?D��![,	"у�N1K�wJw������w�;Ĝ���anR�,�"�#}K6�(_���F,A8��k{U���ҊJ:r�'��'��=ۂ,��!��b�zS9�EN��n���b�=�?���A܍K;�:K�����φM������O�K��Q-�j��
8V�U���]*�� O���ΤXi7c��S7���3�{��`�KdǢ<}a�䒵O�/�D��JDIb>��a]+
����4�ğVl4=��;��Q��Ww�Nf,��l�jz6͖S�c�!-�&����c4��������������Q8�s7�q�}���ʕ2�{�[�,�_�A�f	��6���p��|�uGj|����8�l!��?�jit�G����i�1U݂%�(�y������J�G��9�`45xk.�r�hKO���o�(3IO�Ь�ބ|I��ߐ��mF
	"��Q%K8�rW-:B����c����E\:�9䢣9��y��<�����x�Q�k��?dC{T)���t$g�OnϷQT��f�v���n1�pK�U7U>�w��X��J"�W^���^j��C�?�3"���1)/���v�\�,L#������_~Q}:���q\���)/���?F��uiEm��}fw��N�q����ƀ��zVxd�a�\ov�b��Xq����t��9Qf ���R�9?�����Z��Gea�>���N��*�����T�ڻa�i�����X8:�Z�<U�^p��Fc�=L���Մ);@�\cᲫ�i��d.�������&��)�Hwl���{�p%ia���F��M�����+L�r�z�L�q1]�jj	��n�[`�*�Xʜ�r�:;{�&��|q������y~uN��Lbu����f�����z搾UK��}��k��]Ŏ���ϰj"J\Ez}`�Rπ���<yHR�%{̆���E�!�ef+C�3�$����Ӹa���wځ�JE{Wq�[�\\Ȝ�ŏYo��H���ԗ�����b6!<���I+�?�OH1�m��(����k^>E$�a=k Vl�q͢�4T=1��>��;�;n#@�A�����@~��"Q�7�I�����A�)g���aiY�y���Tn��J{�:�L�%�%�Ť�	Nc�)$���c�ݟ�[�pl\�������vf�u��b���d�y�9B5����j��y?j,�]��n�g�=!b�ЪNIp��ҫ��?y���� �<����@��L�o�yb`�p�	#~��n^�x���g��5i���.�<�MM7�Pw��K��I� ��Z+R���e����5m�R�Hj,>��&*'���&���L�����A�<$,�h"+�J-8�L�6�En����*-�DHU?��&J�B�&��?�X�l�Ij��%�l'��IgQk��m�����jʒ���������Wn3�<�6fG7?�!f��.�3�(�ؓ�ZתYO��8&X�+d�uk,�6v�ƹ�0.��M�1�JGNh&< ڊG'"^�
�wik8N�/t��@z]H��-�CD��I��\���Ш0q�z�5	�L����S��2'���)[u$�r�.Fx���)G=p	4�-�E���o�F�����W+v!n�~��@�-��ِ3�<�'P�<:T3q�S�?��V��v��}5:�%��Z��3���'��3$U(j�k($�=�xV��P��}�Rܩ�$
����S����a ��G6­��9��&iZ�<�V�����L�(�Z:@k����������wzh�S��IAָ��3ܵ�>�AF��3�:Q��e�^���!w��CNC4<��V��R9�~�H����܀�Gnܮ�nC~4q�����Φ���ӓ�Ҙ����s��IV~��܏�z�0$��O���x8���S�-�J��06�]��سQ��y�,w̂���z�c!V�3��*H��v�<'h��du��{Za�ɱ8�Z�WX��
���ުd	[9���=���P��@M�)-���'��fi�VOa�F��L�:@���I�E\��qv7-���(�N�C��6�X@�A&�w%ii��}q�A�*��PZ&ro8�񢴣���2���V�IV���箙�U~Qs[Bl*�+������+��dё����k�:r�l��cG��%�)o@�,ϝ#0})%>���|b�鋍�w�}�arY'�}}*�q��m�u�b��йe����h����7,3&T���ظC���W�zk2�x�\��NW$#�&V<�`�N�oFd�B�y��f7M��� �e��g	��\�dxZ��F�a?����j�Xԡ�".7C���l�0��Q�_w��=��Z
S���s+X�D�4G��(i��O2�w��|޻�����17�dlʶ����$2��6~��ZH�%0h焇����:�~���T΋����/��N�� um�v �z]|���V�3?2�n;X51��������s�;�M�{}n�+7֒#��T��13*���ٍ���ܓ���mO��"Q�~X�XG:�!8����Ɇ��uzX��=�%����l��ާ����Ӄ�3���U��u�:����z{? >���I�U~�3�ꋻ2�	U��Qf麖�`�։V+�j��.�Vj�I�;�2BӋo�D�UT�@�IG�cd��n�OA�4��X�R�#��H�jIU��*A��h
 #���e��Bx���'��p� �c�������2>�a�ja�^��U�	_�K�ȲθU$~).�M�
"�!��
D�3|ӀLt��#I���H�)*~�]��Ol�9���R`on�N�U<��ǿvpV	�w���1~+(��
J�p#�'�n�/ޚ<���䐌�{���/:�� ѿ�wɷ-��jc��Z�����d�!q~�'�ĉ5}.���&o}*���C^� p�_����B�lX�0��b��Fr�bSc�}l�♷U%���i+
���a&!�6�N�2-8�JAQL���iY^�_��E���Wo2����|������.#�E�[�m*8�ֺ.�"v��5�/��	�f~M�\��Zu�1� yD�k��i7�BrT��p���k�m+���%`d%�6}��$׵?����ISO9��d���)�G�svHƵ�B)�{5_���(F�G�Z��V����0<Ӈ��b�X"�� �V!t����M#��3����i�W���^i�{�4��-�����"C|��D7��?{[ �%")v!�=GV,�ƯU��D����Yp�x���X��6�F/�[
&���y������\���Qs{��Y�MW�v����i^�bB� T�$s[8ϖU��&`w7���@q��ʢ����}U������<S3�;�����{xnH)8���sȅk�����i��
u�f������X�哽{0Ѫc��=_�ϬK'l��H��aq�6Py�pSrEg��7��$\i3���|p�cغoH��F�1��K���Մ��u����
\�`�cx�O��o2FY֌LL�<Ck���|��!RE�-���g���b�M�x�w~��(}޿���K-J+=yT+a�	�Uw=f���04*3�I;�Ml5��'�TSF���r�s)\}JI�^�a�6�C���� �"��C���>�K�
�f,e��_��$:	���J3��J.p���}xGa�X"O��SjJ5� ��ڱ���n��Pg��;|<�d���*���I�&z�9��mO��F: ˊO��,��Dʷ�!T����}�o��A�M�I9w�L���� �Ib"h���h4��<�S���&,a��n\m��7��sd� �����h�3��P��Ct
��O��A�R�5x�(��)[̀l1��\�Z�u����gв���cz(�nT��[T�j�)�o� �O�ͳB�w�Ӽ��#�w���C�ޞ [Me??��U# ìq4����rʫl�!�*����p?����5��K5\���y��~���sp$�w�>=h�J�r\+��y�A0����ë�G�2=J����K��@�H�O����-��� m.��XC*�f��Z��<=�L͕��8�.��.����D�E�l���_�ſ/��b�h���"w)8��'��� F�"#��
�t�j��w̭��S{����yGD/IsO��*,&7��'�äz�SOAt	�x1zM�{�C�f����5'���ߞa�e�ǂU|�����68�t�w�);�3�XG#04��@��b��Z����"�F���l��g��i
|�bރ�KU܏�F���@x4g��?q�O�{���M�O�����s������[�6�#�ps~�����: ��Y�8��Y�R��p�5��a'~2�'��"�M��.�5��6UƁ���/�A��I�����v��RTZd�v�4ߑ�����k����.:���A����~73'���0
J�Ӽͱo���"K%+�B�1�Vق?/�G��b6ٛ�(}q¦"a����#!s�n��n V��C����0�j���mo1A���^��$S��i�c�ԡ�/�|��Z#��2v�ML�3�e�  x�/� � 
a9�iH��8�$��<�ߙ 8d��%B�0)�=�2B۴��39�n�<剁�Ry�
�6F]�w�t�t<]:]��|�(Oҏ�I��"���Ɂ�l��LOf�&��,$��irS5p��g����y�B��W�9�y";�����k�_��/ܥ>���b>l3���6��7�Tky��4�g��3��X>
S�M��"������ZS�^틚�֪6��O>]'�G�`3}/��x���	�Yq%�|���kD��%�ҙ[ƨ.�i��hW�ꀸ�'/��\�B�M9%��%w̅��,��9����x؏m�Z��K��5|�d�X�٦�]o�I4��O]��7��&�������N�Ks7���a������2��<ݫ#{��/'�,Bj@�H�h�Ȧ�ܵ�+�N� A��=�	�5ǸhA������1�;�i�]����`?;ް���8I�u�17c�,A�-�o3���#y�˃���3Ay���?�=�M��_pxZ��#lڋN�$Ą-�2��9~���=�x���D�J�4H�+��2B�>#��q�9��<�-G��i�ɮ�R� 9.@/l��^8D�કļ������,/������>�-:�Z7�9xA冔r��D\�D�߫��n:0��en�T4�> �q,m��W��;�x_%c���{q��z�d%�B��Um�����7#�jĚJ"ǭ� ����\!P�J�+н� ��R��(yթ��ֿDSV ��J��
F*�e:���Lű^�!u��%'�>d���~}��� K�_8��(7�o�@zc�/9yd|xU<����f���u��I՞��3��{�*��>�6�5+�Kd�2�����a�B*T�9(K��Q����=�$΂өC�C��
�>o�1�ۈ|������P�q�0s�j���/F�&��NT$�2��f"3X�������<2�� d�P6_4���a@�:�0iw���x�n]IN�]�[�+P��_�	 � >�
p�	q�3�A����"�%����,$�]��F�+J" �M�m$3�����������b�X�����k�Z�І���{�H�=�;iq��v�l7߮�}��l�g��zG��.y܁�Q̢�v��������5�s M`����"��ˇ<����s4$.�����]gZ&��D���=�a���LCK���i��&��>\���fb0>�k���(��j�n���飂}�y�Pw����� sP��|��s-���u8aj
4;�+�{�>>�Z�������Y]gw��E��ON�o�u�̀t�>?V9&_��J��`9�i�i�7�����q���zg�<��!|���ۣDK�X��Ba��g��[Q�5� @�ժ +�Z���>���U��ؓ��/�g�Mo��F�H-T��'7��M����ե�WF���O�)��񒌒?:�OR#�8�԰H��i>IV}�z1�o�dNE�2�|ދ�AJ$��4xi�5��N��[�G�R��R
��uq.�e��4�;�K#]��{F�ۻg)����T3w(�S���HEGR�{����l�7rm��M���.T�s������;J��,ys��n�IKH���R��d�h9��+�f8s��c�t��5��O���mhv���\�%��+U�����������;���c��0��ȕ+�����JK�Θ�N4��a���uuFNAP�[��<�j;�IR脏l�ri�����E���o�Gq$@����ױ��f�!k7�zeo'�9����o Ië�Ἁ9���D�\�~�됄n�P������1|�^Wy�z���Ogx� Pt���2��8�rE�,nZh����F�|ޚ�>XD��|��{���E|�8�容]>ܫ!ot[y�;��ϫC���#tڜ�l���u�3�q"�E�0�2 <߮�Kv(ɮ^���dOYo�w��A|=A�n�_	n����(R��}�~���@�)Y��,4Q�����3�s��9 �;�T�]�V��ډ�g����a�WƠ�1?��'��@q�3�6*�47�-2��8��l^߈uΎ��fE��̗����w���I�ǳ"m4�|��D��Q-IeN1�5J���Z����}]& f�?����'����?�kP�Y��(B�R���{tL]�?IBz/����դe��m�w�R��,i�����c��}�1��SbJ�\�,}%*�_d�m *+��9�7D���]�Q���!���3�Q��Y��<�.��@r��xx`ɋgS=�x�u�_L8N�Y�s]S'R"�-Y��k�#}U��It��U�o1��{<�&���3�҄�D2�	y�?H"�b���=I|��?�4y�¦����:V��	�6u%����p�֙%��U���� S���%�l�c&ϗ�9�Kka�zҙ���Q��w���sr�gZyx��S�,�v׹��xtE����_<C��]�(�V2]�AP�fz�	~�Ez��5�(%��i�ľ�`���7P�������t\ނ��nV�V�lô8�B����L���G����t�ua3�s �wj7/���8�{$��49�h�"E�l�����aG�t䈮ZW7�_�ڃ��2��,���ZO�9!`Xˬ��w��#6Ű �*�&�zOV-.�RWC��	N|�7�b6�!�7������{v+�y���1����t%��©agu�gs��=mB�rQ�(D�o�ġ�
To�D��&%��Խ�Y_�Ci�Qf�3��8�i^KV�g6x�W5�{ �4����|�e�~�O3�XO렷$���o��$L/}s�?��:bG��ڗd�Ws%i��z�����&ą":CU�c-�4i���8������,�@�!�gko�\���}�m�D���"n0�^�;l�t�P�l���s����ZA���`�m��н�������l�L���; �&c���A�� �W�{z4�$G��;�_$��$U�|1��h���&���9W��tܪ8�?�Q�h�NW>��^֤%��{4���[@�^:';f�o�m��X�7_���U� B�$���E
Z�,�s�~Q�p>aq��ľ8���a9�88�f���v:�=��)_?z�G���;0��:�&�Z��@2w�1'��f�c8 �������x�+E��i�+���qc������c�P"� �a��\@�`�������/� �j�;��0uN���1==���0 B�l�3�J)6��fbd��{/�L�2��CL�l�)��*��F��ҔN����J.�;���D���_,���@	x�I|��dtp��.��ʅ�no���_���+�Y]ʛ����R�]��O!�pYJf����,�CeB#�D�C^��*j�8�9�\^=(��K�ma"Bf�ݦ[�t2��}~P��kGd�!�C��&,n¾�Q�y��� d��h�*d�O��狣����,���V��SZ�,~�
�z��A�B��2rE���n^�"K��M&B౗���s�@���̿ש�ȍ4�Fx��>3¯�r��*-�M�u�.PH�ͻFy�;���,xd]Ⱦ� ������
��Sk RQ�A�MJi���W@�MGV�z/��.�ݷ�uM�$)gR�gUI܄n��ދL>_�x^Fe��f�U��)N�᲼��30څ-��%�̟��͒s�z���H�_��2 ���%����Ͼ?��d�OG�m�l�~���ٗ	���R�����J��ҽ�ܤ�������Lk_��N���2K��od]p7ȱ�EX���/��h6xIs�vL�a�͵?΢3����,�1���#�)���l�-n:�ch�s+*-�m���-_g2pa-�{Ak��
�@��w�d$k�~���D�E1.ʱ�Kܭ�2�rΣ�I�/\�+�d�f=@)4�]1���*8Ȗ�ݛ��WfN�����M'�nw?Z�x�x<�|G|L�ą���ŵ�5�X�G�2ycm;o��uXbPZy	J����E���I9���hW@Tk)I��9a��M����X��P-s��en���h�����̏��zn{��baO���ۑx��\S�|v�I2藻���������%x�̑Kv���H%R�!=|�_���RgS�e��30 �'j�n�Eզ�������U��C�� ��6[T��O��Ɠ�\������+�x�,�(���>=�k��kp ��T��7�N"��\�]f�'�u�t5W5ժ��Ό�5a���:�Pۯq~i�-��ɡ-��H� $�Nl$�Э��
�8.��!3CE��FD_oJ��d�=�4d����z�Ŗ�d��Y ,/l�����1} �X�" �Ӽ��`x�N�8���6K���`1��->]�
�Q�{/�J�)ر�%��t�D��4��L�s�9	x	�;u�a1Ѣ�b4��� ��C�P?�e��!h�ip�rZa<q�6W�D��Y��)�}'��{�k�<��궇⏹6���Z�Y���<.�q�����Ԛ.k�~pw�)�n�B���8Ȧ�0�7?1(-��Mb
F��.��O[Y��[,��
��Ҿs����<Z�+�~��:��%�)T�Ɛ��L��/qPB؁&-�s���x���'k�e9�
9�q�2ݸ���tO������˺��};$|zy�U棟�W�R��j)x��e�m<-��h�
����9�ބ����L��+�n�UP����������¸�H-KD\�N��/W�٠xj�!���kΏ�⇉-.���'�f��>6�OoSU6_Z34o���K�rPR0��^���R����קR;#�S/�!>]\��T;����Ȋ��m!�鷬�����*:��0�U�iI��0c�~�B�h����aIG�Y�H�=gp�xC�61'���@��:v)�����P*Rz�ٷ��b�n�y���48H��8�]�Pf�Rj�`W9YrP�`���)ɥ	�c�)��:�ޕ��[�7x�*M@d�e�^g��c�s�u�7�nJdpA㐫��)��м?R����y�����2��14MX����h�޽���q�_���0$ݠTbsz�'q���#��;�k��m;h��%Ug/��������o�M���׈����rv^w�!���=\7)�����'(�v)��P�S���f�������A��.�RG/��,��"�dQ0o���f�#(�{�:6E̩�`60��ND�}33��Np���F���`ۧg���j��&q!Q����L�>l-7�����F��7�řJH��l�O�5�����P��_�_R�����P�O����
*��̀�
��L����^Lo����1K�f&�B��'=t����a^���t���qo2=���@=r�B+�2��N<Tr�p=Цo�'�Aƞ�,�Lx�or6�N0�f٣�h�nԣ���f�㖢|OZ D���O���bA��828*�Pe�������@��e˵Jk��ȥ#j)N�͹@`���� {k��غ�`������2:�omt�e�xP,�L�������%ܡ�+�4�'Z&�uY��C(��3A4ӗ�d�}�Yd�\V�.ƣ�:���ėDgޞp;��߲�_��ش�@}������)����&ۻ���Ů&茉��fz�T�����I������U�X|I6#�-�\zPԊ���2
��8\v�n�Q���3���~�]:��Dnv��.I}b�L*j�j��٭/
y�YF�i�,ȳS�N�S������,ז�v;H6���U�#Y�;9wpN�r#P�CY��n���_�3N�U��������q�	���"��{����!!�/m�=�|'k���*JP��ﱘ�7��$窝�c���Z�#2{t�SN*���D��}) �!�$�4�i��T��5���\m��?k��2�$�2ő�NO�$�eQ�*�:��4�r���I{}.$ѷ�q�)/���wĀU��v��^�n�����R?�㟥)�g��B�ߗQ&l��#��4|в�UY�Z0	��.+.~P�<5�*��f�ЎRI��$�A�"�T�.�z�D��  ���$5�y�:r��p=h�}���Kmpa���~��j���e�ۏM���ծ1S�K�X��8b1I/��`�vzD3��!a5F��v��N�v����y~��j>��)�xU�<Mǝ�)�,+�UV��.��$T2���W�.Wn�SE�&b �<f4��j�d���h�|x�d��`���U�~�{�?�����6Q&����!��O�w5!i��P�ecJ_��E��i'��})e��2Jb�#����.�?(����[��sW���(�ᛎ�o1��^����G��ݒ�}�vó	��ǔ�J�rȽ?��n���jێ�?Ka<���s_U�L�H��{��п�o�Ph.9��F���	��CfX%5�)/c�J�9�"��KkH3����?J��O�eQ w:5���\��
;a�f�S5�3����M����$�ɞ g� Bշ�M�F�#�'&Ƭj?���(��"��$�htH%�Hu��~�h9k�%2 E�(��9W久�M���o�r�A��I4�+J9���Q����u�;�����%圡�q�Uós�Xr6:G���bo����D���j�n�Ե� ��p���8UrM
Z�},��a�
���C�� �ˋ�L`2K��r��	�� ���872Q3�3�D,����z"2l6 CN$�x�Q�`4��C�� K�����b�AwF(g����|�^�f#�D`��dF-[Y�n�zF'��}0�gԳ��ph;��lg�¦�e�)�w�V�رv(��l�r]�>��M����zz��u�_�������R�*��n���0��w���xl]8a�3mG��y�zEn� _R[��r��^ĉ�Oe���a�o�B�,x��ƒ����\�k<�y3|�s@�J��+�]�*�"����l*x��~w����[�n���X���u�}�
ZX`t#��<�.�u�)�>�{kE{2w�.�d�k��[�.H�/��%z�$H?���V��$)��P���Q8��Su�m�]�_~�7t럡�!�T���|�CQ�e�xpg�Ial���gᛨ�27��9�0����C �������;���9p�^�ۿ�E�*fl���o�A&�h��EI��L�i�Ж���x�Y�ʀ���vJ3N��7a���Տ��d�n@��[��A�K��H����\�&N��oF��(ړ�Q�Ɇ���l�)�Z�Љ.��2�u�E[��r��.�S�D{]D��+��q�/��L%���l��а�D�}��������3��NF>^�M=����V?����IH�\��z ��=)��,4�F,�{��{��g���7������\,T �4�%�Ƈ4��yy����76?f��>�O�.�m�T_�H�����Ę���C�{��~p�T�&Ƒ�6��=�ɟN��0�R���2�K��t��1U� �'�]��|�܋�:��tF*�.�q�LT�_�h�F��:�inmY�����҄�o�fQ�2^.��B�·`��S����1����h�f:&\?�&�"�T�R�f3 8�/��"rx�[M�>�����m������/Y�����a֙�d���7K9{2������FV'If�Em��sv���?[X�����GUB�𺑖�Ϲ��m$3;H��w�{�\�Z@YT��>��A�I01rDyb<���A;���(jA�;�v'��Iު��Ψ���"���F�.�k�\ƨp8u��u`;�AT8>-�Ǟwk;!��_���L����Zz��!�n�cO�I��X-3ͺLg�)��;����ϒu {NT����%n�f�#ٛ�t/��{�CP��Q�"2�oq�ļJ�Zn|��B�T�PyBQn�XG���=vR�?�c}�� �tY��2a����/�
�m�/M��c�?)%�_c_��vG���,Ĝ!���5ք��l�ZEؠ����T��U֘��	�&��2����=����a�(��۪'�V28��\�?,�����,(
����>b���
h$�#�+'D��,VϞ�"m�AT���� ���)�% o��7�ZC��_��M�v�;"�$��疚�F�ni�(q��6?�O�8�(�hT�ʾ��"]�I5(>zmq �g�d�s��ߋ7ex'���A�� �u�zoGgq���ͩ|�Y��k���鐔���/����el���mw����ޠH�I�Ew�:l����jб�l"���.'q ��À�-Ӳ�R�	���3�i�b�n�%Z	�?�%G�=�`"��$�[h�ſ����	t����՛I�,J����ov�7zB�]�V�o~�o��X�9�6�����t0�d2`yy0����%(#%8�(��S9<���b����z��,�L�Q��W�,�)�E]8�3}�]�wi�n�@������|΍t?�5̨#�/��X��$RyE��[�S�H���wV���M�%[k�<��%�>f�(
ZZv��w��'*�l�M��a�}��Sj{��!����[�sA_W���lMZI9KU�#B+xS�T�צ�O�TNF4�p���� �{��g6���3�=J4��%'$+�J���]��mm�am�uWD�6�vG�VP�U;�j�QS��l��rI��i�OfJ��a^-�R~�6!uɖ�6/�+��Xu/��7� ��}L�<=d�`��K�^���3���B�ŔY����>��E>��7�������'����� ޔ܌�_�@����^��!(i>[����p�^t��:䵓õ�Upf�^ƺg�q�J	� ���FJOKb󚐅�p_@`��ט�\Wpd�g�|���x�0S*�� $��:��1���!��V��xtƢ�Q�#_�������C��~R������ǳ��z���ë�PN��l)Z����n� �ɺQ�W�.�&v9n�7
qa��W�����r\GPo�n:Ew��=cZU�5�\Oᇷ.�!�E��0�>^�v��F��T�'�$]�5�+�[���b^r#@A1��x�:2�#;]X�}kh��d����[�;�ܟ�[���⹘���P�v�F�˓f�m�X8��x�c����NPR#�.�[�0��H��u��ng:��W�h~tG����W?��1�V�$^��1��N�	�\</uw��F�g���nY)ƎYsm�[H���~�X����P�\��/tYv��p�i�������#�>U`@;@'�"�\rW;�D�L�0㳍Q�/I�V:�b6駨�b�*��!ێ5kw*�fE�V�\�ͲcGX&��R�\��v^��`[����F?�����m�!�.�br���oS��P��!j5<��dN������v�o�`d���];����!X۱��8 y�6���Wm��TI]�[��n�k�A#|�[F���U���A�e�?{�5��țw�E�J��""D>bl�W8=İ�'�Bw^	4�PG���%7.C��#JڑQ#���0�e8�y����w��Z��w9R�`+5�})��Q�N���ΉA�������2�Ad�]�BȘ<	��"v_zt�����#k��rK�^"7 ��/�F߸���	sl�G:�B��D۟�N>)�|���+��Q?�E�X����̪�"���xoD�$:����;�Mر�������L��}o��t{�q�+T��P":[(��O���2��ː�/i�Ͷd�vkݫ�x�~Y�KW��i��F�m����.��ztZ�b������{O�����֞U�D?�vg�ؽ��^$���O�04V�%-F�:��k��j�<��0ፊ_ޞ����oZ{��91���ft�^��o)$��5>�s2��������"s���a���/��6p����T"��	�`�<��6�잆�r:ԥ������e�Xv?)�E^)�hg\}ʃ%�תPQI�l$O�W<�'�øk��>l�o����wm5K����eT��X���2@eV�	c��%�cN��H5��<G2J^�w�<��B�y %f��K��"E�MX�R��$H܄͒E�>�#����!���޺t�\ �Ca�䖗/����w}c+Dx}�J�ӣP?�!O��Zx���G�B�e���E=��i7V�Y9R|�G����Ӯ�{*��`P���_�v-�5(��>��,���7b����d0�:��bJ+���a�*��ǚ0_��0	ɷu�BU4�����5@G:#�����L� k�m��N��x�ߥ����Aľ#�}w��E�j�U�
�o����
�����ri����pUAE?ģ��6�3��K��U��i��o"�G_��x�R���N�GF�@qmuFZ�,8,�j�s0n�qឝ �c��È���=�V,�i�,����%��q
t��H*!��h҄K��~���$N�D��j�NT��LxFp<�å�XOk�bu/; ���:[�j���;��|]��f(�0X� _���):/�~�i����Tv�<=�,��&5&��\loW�NRP'X���������ZL��i������Q��:ԝ�OqQA��GH� q蚐����_�6����3�@	���BR�zX<��$��@�6��^O'����%@;t/:;���o�h��[L- ��!�&&$Ԏ��]jD�|M9��N��g�)�C!��Ux��N�5�%on(5���G�"��*���΢cn�8vq|O���D�k������gA)m��+����Q�g�个��X�c�E�S	�];��_���aQo��XR�L�5�{�+l�����bF��=�r3ZQ0��~�[8Ȇ�����ܷ�PW��Rٜ͠�0?wE���]J4�u#�^�۔[�H�37��=42O����ۗ� �&ӗs�U������9��6z��;	]���D�'!���x�-ě��� O>��3�����A��a%|�]������}F��7�I������e��Co=��:�Ϳ���s�$V9�p�IJ���W�b��c)�����FU��-����Llo1��*��9,GL�@yX8���ӣ����6�S��:���<�*���K��/���TU�b�)�/��X�����p!�{�N*�S�m�q;s�]�5/����c����(��h��F�;̵��Uʆ�?.~��������*��	Z���>��6�~U2i5��;$��<&� W�#�c��ƶ�"4�S Z����k�ca*9��mּ���>���Tsf;8q� �|��eT���%䴎9c�w�`M@�
h7���`�s_L��h�J��/����5�bz0R*��T��t�߫ÉqҺB���R�a���E�����ըMa��}�B��fH�e�z<y�,�jr;l��&�\����g�pXBk�� 5vS���H�f���R.��d.D�+���y�3]N����bY���[���@���>.e�g���|3�&e�m�B$�>�������-��2{� O�<�$�E[u#�B��T�W�6��I���TD�=GM�moG���d+?�_�(	�3ju��ߊ��%G���=�TP��:eLc G�7r<4l]�&Y��/#�e񣿺
mE�U+<»W*��5&٧��o�On�N�Rq:Y����y������3z}��Ŋ��{�X�]++����}�9f�yLh7Z��ɱ>����ָeH�<�-7b�G�=��Xq1����`�E�4���Cգ�2���"����pV���ة�(	�]�<���*�		�b��-��Д���$���Qbs;,Ķ2�X�j[�M���������*faQ)��g��ݸ� To�0Y���J����N%���vW�|ʉ44�ݿq\��������F�`��B�iMG�(J�J}x{!	���"Z�!q!co(�y�
���+�,�� ��0���K9u�e;�����%�jA�Vk����vh�NE?����B��<��C��ѭ����N��3�	�m��{l�	�_�k;��U�-�c���ǽ�9�.�c���4��4w�<m�sI��6۩y���k��I�:�������� �M�j���7;P�j����Oj��DU�6B����#3�$5V{Hh-rܩB�I����ok(n���Lw���A�Ő�g$mS%�?�ʲ�"e��N���*��l#}[p�r k��"�W6C��:ȿ�ɶ+�:�2�K<`���U��z�'��u��6�����!<]�s�%~���T�ôG�=�=����*bhkʙ��"�>�5K��Y�l&��Q5m�Ws���'m�z��O�0���)p� ��.6�)�0U ��L9�65$}:WoX���葰:K^��B�#zB&b�_V�S'�<��DؗbL���+�㎙���d"��d�a����r�_�������<�$����P,f����3`�О�O�i|�H�ŧ�޶������+S�;��a��5��������	�ڍyE��"�i�	<(��.P|���¬����7 k��؍��x�H��������)J��`O��<����?ԧ}�c�8͆�����,C�ڨ�|�@(6@��<�ՄǑ�;��A 23�OG<U����t��$���i�!?���}�������+�ѕ�<'4\�����L�g�<�[�Ud>�,҅��3�v���B>8}o&����qH�g�/sr��l�6]�����U�&�aר��*=�*�~��8B1��<W�O��X:c�5�X<w���.��f�hx��*/���j����b{�č��,*���'��j�:�6��V��o�����v�'��?�~Z�vA��	^S�^+�k-��˧�<Ƹa�PGQ.T6��0E_�{�$@Q�� ����q���d�������HB�<I��IJ��ze��&*�KITKn����$�lq��T9�)�����h�LQ ��F�t&��_˟��f�#�Dd�a	�N+K�3Xq�X<)�~��:����1A�����eʧ�����;�ʘ�����v��3`T���5����@ ��.��|U����DviVd��/��{ژp��+��)k��zo��7����D�)�{UD�8��$x�Qg����nN�m
��N5N��I����ڀnlB=�nO{��}�<|&���>3�CM[Gr>Vj��BԲ��,��e�6=�C+�?��$��R����_���AD��q@�&�T�yS��W�k����o�}��B��l>4L2b����%�w>Q�~�vw�BH>��"��Mw��DGDW�H(��!�/$+����o�V��r�VRrn䄻�lZ�ᱴ(=�b�_�m���"�����+}�#_�Uq;c/LH�[)$��qs]7u ](͔�o���5���u���KrȈ6Gn~)G�/4I��BPf�]t�
}��}�
~��1l�<�%X�������Bk��D�F���?��dJ�+V���rtA݁�v����G,��x�܊�A�I�i����\E9Y�}�FI���y��L:i ��_��	�V�$8��jя�W���	�����r�^�u��c�6x�`@��W4�y	�[�^v�`T��c����x��v ь�nQa�l���z���tMi����1���.>�F��v>ھ��<ոAH]� ���[��g1��"�E:9M�qI{�,͘�i�/6���u���aG���η���ޤ�i����6���5��U��pAp�Z�gV�u��>�^+
�s9�$lLi���w8*�ᑍ�iܠT	�KD��s�t�K�ܚUXK�5��O99��.����;����Lb;�ͦ�pOƮۭI·@>�`�5���-�� �ZW aýGz�2��j9p(�V�ؤcu�c�]�Kr�Yɓn	����x7����V�j����	z��N%[[/���ɓϊ ̷G3�^%�J%��N�5��p&�i�5`)�?3� &��]����W:Ө��OJ׹i�ƺ�P��I��W@K��/
��Ǒ~���}A>m��N*��K���C�J��iܤD��!�iֈ��f��������	�L�;J�3�9�m�W��Z0(��,}���(L??�*.7|����O�l3ȏ $O�'�a�<�Ƈ!�]��:ضg2V{$6K��P���ӌ��)3#aO�JgL)Rc��E��-+ƾvG+Ƈ�L:�5^�X�^}m�;�#�-�	N��A�6�rX��+��M�ciڅ�f}=��1�8X�������9�ֵ>@,�����$zB��Mλ�O�G�P��3�4��!�ڷ"(��Z��T��Đ�]i��%^�Ȼk��B�Xݾ���>�~/C�U�{8����H�z�<������E��im��.�ؓ��̚�@��M�|dZ��
ڤ~J� ��&�B��)�2j"����N������4-���[�v�o�>e*�.r$�s� W�9I?��bZ1�ڲ!u�F/O�i>�r��Z�
P���j=P뙽�wd�K��,���P��\���2S}%�
-Z��0|����8�8�L-��pd���ީ_c���8
k ۏY�����@�14$�v��Y���J��s�W�Y��sSF5���s�4b�F�Sv�ͳ\���� �{C��׮go��\3JK�*����y4N�
��A�Ji4��Dl�@�|"�]X�,�xa��b�V8����㗈^ߝ��)`3�e5�)n�e5��&�,֎4�a�P�G��0�-�<Rh�2gy���9S�հwv�Q�s�W�W\�vk`���Q^B<*²G�mC[�ݪ T�x��J��d�Fse��j @��Tk�P$� ꉯ�U:+	�7�N:/;����MX��/z7)c�D�9�Yls��|�}���Ԕ\-כ�-��=�����%�]$�[i@�E���M��Q;���2C|�P��,N5�
�
�.3�����\N�j<
v���E���JDʑZKb��;���9&À�\^����dbK����.��W����kc'�s��K�r:M�����f'�����!8*�2�K9�o�| vxOZTΎ���Ŏ�~4��*G�ȧ�I^�z}�����0���t�Q��３�%`ն�!f�~��$4
y�Ze,X��t�S�H�;�օ��v`�q���U�n����K��E�R
�b�y��wcH܇'p�Ϫ�ڈ���7Q�(#�`�"�%ZN��[V^���25�/�߳I]'�@o�cv��I�
�ؘ#����Ae�����i;n�vA>�p��(;�p������V�-������G.b��e����~5E>��oLA�|Z����i

<��_�/o�+��U��4_kH��n��ŭ�K��ԏ�l�J�:!��C���.(����a��lX��`s6�H���cw�.j���K^
i��Fe�%Y���%(py�G��q��쏎q��_������k��P�?��T�\��IwV��)n�^
�������of\�O�S��_[Cp�2�*��ls�0b(�,ڐ��ʌ���5ur�x�41
W�TC����$a�|�hM�~$<,�=&�f�Z�����A ё
��о���E�O���i��iq ],8~���\M�E�8�����Hq!_c�D�ok��݉�l��լ:)PSA��b�
a��C��N��B<�r�~p�:��"o{&��R�/V@Lo.@
�|�-��ի̣�ˀ�I����F����'�Xe�ǡ��(�)Q$���	2�?�&ח���~���J���/�2��5�23U$P�ή�Q�u$D+6�Y$gi�G�f@��}��<��D4і��_���(� �Y/TKOE�Z�X�R��?�;�na�
�m��Ȃ{48�tMk�� @%<Az�X�e�B�tK�E�7g�?��Ԃ��~:p{|V<��k~f�o@k�w�BdE�=N���v��'%|�ٵ��_��h��`mԯNS�'Xu�P����1nKi�7�98h���i��R�,K���w�D&��2Ri�vs��aw����9�w�1�m�������Й�.��W�A})�.�Pt��;y�0��կ*�/S�A�k@���䈊�eu���4s����;��C��N
��J<�r?���f����l��6'�~u��(!���|JD~�V�e��*���l��8>�.���t	J.zRg�w�P�e��U�Z�Jj��Щx���z�M0��#G�L:���^���?�Ewp@z�I{�d�g�^�Q{�2�����^
��Q!.�5�\ i_�'붘~��ՠ�Wb9�ʣ��[j2^��'q����X^���@ۘe�y�Ӭ�Ůy��3���NO��vu����HJ�Hn���z��w�jbo�-.Ya6�~R|8Z�
VE"��Ypz+v%vm���
^�_�-I.�قN=s9�!��>^c��t5cG%O�G�O��7����ID���	؝H��SB"�ΰ��=�m�L��U�^��w��L7 1�
P���05e㋜ewس5�CI8�㫄���D����C�mH�ެ 3Ӗ0F����iS�s�-����6��\綤�������u��̀G
����_rNu�|k�sV������n�_���t.�3q�E,n�G�k�E��&���nbm�Q�|��}@�/�Φ�ظ��Mp5	��{���Q7�9W5�QjY��;�"/&�&���y�o�- òG�|�ޟ`���c�����Рq�k��a���G_-���-L�:Q�j+2��� X�� W��ryv{n6�>膵<(����еk�z�������7�DXw���<���������Ϛ:{gvm���P%t	�?'V;+�Xu�Vd_f�XfK��*�p�)\[�Ц��j���u�u��T��t�b�
����9@��}�V���Dw����j��N�I���b8Ov;ą�Z���X謹�����M���ӈ�/��\n���5@{	샙�М�����2�Tؘ�Xؑ*]��|;��yEC�#<3����*���I��9+��[�:�t��@��P�Qq��\��}$�ֲ��,yk�.\l7	�z����w���<������!�#2�C��b\���T��\�����������vh�Y�-Ƅ���H����ؑ{|��@����+'��� ���dLr���7T�$�>/@��~O$u:v;2���*����Q��bDURX��4j��v*��m�:��\VO�1_�z%*�B�koM�a:fK�����C����}>f�����T3[ݙɏ�Y�a(j`@�@\�N�pÚ� "S�B��a���� ;`�sc˟�5<�\�0�=+b��Ԟ�	G�� -J!�0�{�W�qbv%2/�р��e �('ã����*���v� D���4`��=,�e���?81`���X/͎\g�플h�Ղp�_.QI�HY��{������eb�5_���A���ך4$3K������Ƹ�"����X<>QD٨[1����9�>�W�o�^���Żiʐ�Aw~E�ޠt�s���]Oh��{b,�v��U�{���.�
.N��v�
��t�����7_l���bd;Ws�r�(��BN�vBɏ�Wi��i޺�����G漐��:�[Fo��r����	%� ��3R]��Y8pƬ�Q�,EM�U��#����K����̡|�$�/�P��%�� ���<�i(���!��``6�f˶�vC�y�����3�Ư�^ ��v�{��n�TT��8ǀ��Y��y{��'+��)��t��eT��Y|i�{r��b}͝�<��]���-��Hi�%^TXj�'rS<���h��.��i3nnR���ì8|����9�f�Ⱦ޵A"!�1�x�)�=H�v<[�#m웉�!-�"G�
c��Ѹ�U��7�R��	�,p�HG�Og�L�D�P�*�!@w�5��m�4�I�5�t.ϲٕ'8t���=?�ޖ�Hz��(�W�V�G��U��Vj���Wn\��R�؞{t7˞BO�̇�LI��ĊOBX�%��g��1q:�)�8Mn��w��%��	�Q�؎���<K�EQ��� A��Bx$1F�B�r�Pq��f�"/�z��
a�	|@�="���5D^'���ҥ������D��+����֟�О�pWn~��Yp�F�AhM-��X+⥆�L>=S�`�܇�Oչk|H�f�x[o��U��=P�]��d�H�Q��a�&�H;ɥo��ꁅ��wJ��u�x)ͅ���7��I_ͬ�W���f����m���H۱cӢfc�6���XI�&3d3^ױ�/�d�O�{��#g�����ɢYb���eS��+R��A�ޓ��KB�M�����58ѽ�����:�`�D���]��P<*�3�AB�Y��C.��Dô�~��I�d�w�x���#�:=�̧�*���80l� U�f�	$����8��2�R�J��Y���oT��'����h��E]�o�Z�`yǊ5�]��'L)S���n-%�����y��I��L�6(qp��?z�_F��qV܉��\����Uf�j�S�r��|���޿f��D���\�X��p�P�R3�R�v�0�ms�D'��7���7��@��F^К �K��:u	هV�7�G�
���Ј%KC��ߢP���U��k�Z��l4k�ONGU���I3tڶz&�Y�4	�OIYk9��9���n��W���3��.JX�\���u���H���!�jR+��|�pxt����v�8J�J{�	�1syQotʌϕο<	�b�l�và���yPc�,��xA1�~
b��мE���A.�^O���^�d�Z�ۙ�h�0r ݙu��=�i54Ӝ3�~T�"��Ti2Ͷ��/�?��<��C���B���v��c.E+�ȑ����ؕ��ˤ��/��z4G\�4�;�tHq�e�F�R�A@n��δn.cnKA�8n	݇����G�t_��h6��H\�fQ@]��Iz��W� �~��OS���F�e�Zؐ1��Z�l �ޕ�Z
�Z+�3���D�����
]pD'*���-#��n��4��!�w�,����D�<��t�P�7����d�I޸.�1�RJ 4N�5����ؤn@v�ڰ�qc<mYZ����䆊HN��D�����%�ڭ�r.S�����Z!����{��kZǷ��j���Ն6�m�؏���^�.�_):��q��V�H�H)R���4�f�H/i��k�u�b�N'(٧�\GؘE}�/R:+��-P82��Ρx����&ʺU��șN�X#.����z�����BNNx+�#Ǯ���%��"���P���J5�c��7��)v�x��������F�h���%��P:��-�c�;`�E-K\��e�6]�}�F��ɋ�dsb����?��!F�*��U!U������Wu��	���Kw�-�L�N�n�g�Q�7$�e�j�*'���e�@��V���G�֠,zw�.a� ����`t�'�	�Q�Q-h����`�^g �[�Ƒ{���n�'ZO(&���43^�Q�/�rA�;OBC���H�I�"���_�烴O��Aw|��4��Ǧ��Q�q�Z���dh}zz�����M�^NBW�4����b��gr뇌�	�>�s൫�}eϦN�^���XF�a�'�[3#�fs��=�?T#��)?G N%r"ֆ���=DFM*�+K=��CQT��;)+���\�F��l�?��2�z�j)sg,�kۆZ_CFU���t�Y�4U(YݠO����QWFd?Q�� ��S�J����S�,�6�"�=�R�`nD��(1:���-�+��! ��q�\d�F�	��&�{��?g��|��.1x��Sl:��nb�"xZ��-�9Oa=�77����T�m ����ItBsBG�^U�N��q^����\A���>��]BRyt�,���R�
�f6~2�b��΀"J%��� �W؝�d��ڪ�s���	o��uKocƹ�@5۸��R|'B��pd�����O���C�3����;��w�S�uL/��w#�{ϛ�+�T�(@a�1]w�Ө�fJn���@��;�zU�>ܷ�E"1+M�Ahtj��_m�AU�_�>q5��L�����ʝ���e���C��Β�������y�H�&vbN�Q�:Z�6@��C�l�*�荆,"�K�x�/ơݣnY�q��A�*�¹���~=������rRv�r���H4�n~�NAB��ԓc�Z�R�;�el�	$���!���袲�D�/��UK�0�_q�^	H{�I��IɃ�����Ƹ� �[� ��wu��F�i��bCr7���|3�`�I��y}���_�TpHJV�g��"�p�D�-S�y�vM�)V�ZG�è`S��BX�d�@��O�C�b��;���P�d��G�$�F=
A;�G��|7�|p��.��O��$ �D��f5CӃ&KMz�;ވ-�� ��iko��Q�W��O��-춅<�&x2�E�A�"�\C�`8{��x�2�{�}YT0�)���x���� �w84�s+RB�X���2���~}��-�)���8yz4o>���I�vM zr3ʥtӉ�|��q�^W�̋z�H��$�һjE
Y_lh���R��kar�6����Q��3+���q�U�o}�Ү�9&���-B�C�I#� ��çr'�0��Ʀ�4��Py?���ja�����Gl.�%t�D!�8�)I������B�E�<�ьjh?η�؝|3�B����j�&.Rin��o[3��Z�����ʲB�� �l3��NI�}�;��ײ�F�fn�w�����?��G�,���"�ŗ?�_��w�_�e� *38�mg^'
~u�p����vj'�<	Q5�@����#�H|O�	�õ����s�!*�'ɶ÷z�0]��,�K�� b���q�h�\�A_ �(���t/��p&��h@:-�G�rݮ��]P3��i���F���m�V��+�
얫u��vV����&�p�5�oԣ�6���@:OHv��!�I)�X+���g�(ے�R9I8�Gjj�euX��y�)i�x��bd�NU�|8a����b^ǈH�Q��i:^4="���v�����#�}褣��H�D�]�q��K��0d��z����m���2(�w�~܉qP�OTX�cVe��U�Ń�%��X��;�մIeh�`�(�G�l���[1{7�Z;�s+����dq�����&��ߢ,О]�Q�c���
�w#���[_%�w(I#-C6��q�<9&3�s��k�,�GSva�#MUZ �#G��J3j�gN���j*6����&�ޡ���6v�$����)�v�<���q���P�����.(�ɏ�T������x�cn#�<�w� ��w�Њ� �{�ص�s�8$�=��HU�=?F�x�UQ.�w0^��G=)�b�Ƚ��KZI�~������)&3�۽���˝/�l��������}Ka�Q�������׾GG̟�:}���Ư��}����.�h->*���>`k�hݲ�s�W�rE��)=0DH�/��7ݢ����V�Y����M�����xN�k����Og~���F���Df��3��{�j����D�g�$2	��Y(Ù�&&/�_�ȗ?
6�5��դ�H��sS�&�|�����r���Gk\?Yg/�N&������<:1�j��"�=��lF>�q�O���<������ʟ~�MA��;�B����S3�Jn(�T��Ȯ��LFB������2�4���@1vJ�����~*y�d����i�k���ij��	�j`�&����G��L��W��xƬ��Ϊ�r̆�XXqrW�<W{�Ğ���"��0QS���~��Ơ�0��0�㺥�V_�o��]��oipܯ������/�a�v&EI����@ߋќ{8@�������{t�B��_�3X�����������;-lP�i7�M�T$�S|
6Y
.GH���U��%�@mn?�<oe.�!ZL1O��3Bp(n��Ae�Y=������LS^!�<�_��Ҁ��P�A��/ z*��; ƿ�K�D�q��KlH���.���µr��!��~ƕv����mּ�<����O��f���b�:�	���E��5$>��j��.ot��E�̹�!2�u���UZ�F�����I������|�o/R�Q�8�4V�ۀ��݇�,G�1��)V���d�߷yP�,�gپ=U�݆T
�|�_�p-��=ZƏ���-�&�}m��b�V�["�R�)At�UB+}X�\�`�Rz`�׃�jW�����)��@�F��V�S���'��7���K�=�8�HOGQ���Q�8�2���
����|gla�B=@�y�����w�k���wɉ\�Oiy'�A5�g��:��&�̟З)�<t�!��C�غ�q3Ҋ��ť��Gl4�t፣�R5��~��m�ͼ���sW�{?0��eԗR�u����0�7�����[�s ���8��_����8�]C��$���k�� rG��Ps���)�`_�"�oM�,�!�3�֖k	��s�P}E�
rw).KQ���M���I��b��M'�7[�Y��=~��{Q���E�~��ϯt��t��v��3Bɚ{d[��'ş�A�;�M_�֜�s.v*��O$mq�{>�t�s�B-��n�\2G�h�z�lj��<�9aQ�1��bJ��}L���@��'/Hz^4���3�|�V�[�k�H�xSg��-�|}��8$�WƵb�4n"�w����R�4�$�_́O~
۔m��h8�L^�Wu�W������V3�
N�l�S�=/�t��cJ[��A�V-��뽿8ձ�#hk5�2�00:�`)�ifg7��	�ȭ� ̀;k��_��[��VտP�	��B��h�ˇ�����W�gIL){�R�4��9�F�(p�F�5�1���uO �P8I%�U8��ވ�ki�� ��W,H>v�@h��M'i8�{*g��������@�j��R�8���q��>i����
\����~�(x�7�x��ݑ�0�`ce��b>�6'�\zd�e�`%û-xNai[�B+�6��z�ɱ��w���9�GOˆ��T͟�)�d0���言g�����t=��*�'L��{=))�yo�oS�
 Q.��0Hҍp�^���X:u X��̡f�����?�=L�����d
��h3k�E]|1� X��X3 {nx�Օű�ɗ�C�F��sy~��f/��/w��C�H�������s�N�s~�F`���*9 8�^��y�0s�4Z�b%\_���x���"��"�
x=Y��KUw�BfS����E�J7�|y�b(����i&����~m�ax�8��!���j֖�'䡵V��'���&�h����:�F��dQ1$Vg��Ӕ�wF9w���x���N�P`��U�jB2�ٿډ����
�ۜ-�bNI*�2�*�Ս�,��nR,s�C@�1㡴�
��H�s���@J���̃+;�ޑz�$tY/�ގ��wU"���4����Q��p����k�{�^xx�I5KB��-H#-�"�jS��l�o)@�q�m���ߒ���:+��r�gdZ�$ks��GE�1�4���r������ ������K*W9�Tm���m�
���u��?��*w�(sY�P2�h�s�D�A��j�,�L�o~kՈ1�k=,ѷ�p��IT%0ҙ*�����z��82ن��p��������$�4�!l��>#	��%^�Rԯ*�'�b�����[�f�C˫zBv����.Y�ٽ��&�~��{��~�pqw55�J��d��&�=�q!m2�;�I�KS��:��>����$ߡ���{e�n�u���=��z���$f��7lÏ2E"�0MZeC"�ydFo��.�Os��a��ʯ|u��1��d��f�N)�S�b�f!J;ZD�����e]�H^PS�\�(6��}/�$�ٶYضV<�3|�X����_�
��p ��܈@Dz�k�x�AS �($Q|��}�
��O	����%���X1���Q�p|���[5r��㔦��7&"��|����xZ��O�Fղ�;c�+�eq]�J���w$�4Y_A�s|��S��ۢ�3��7�P���3�3
�|85{�p�A����R�S 3´=��������wM9�)b�F/���T,���f���g���	ޝ)�7�L*�#�^���� Uٹ¦܄��g!��'�T��{q�n��l���7��S��Y�9�?�Ӑ�Xv�e�;Q�d�UO�ˮW�x(������Xj.�1{.=@�`�<�I�`�K&?<S��ʒ߲��gx[ɷ��]�E!x@�]�,u���6F�;�0y.1[}�߄����\���-�����ߞ*���;�]̩�����˿�K;��޻�m���Ö�°[����H�\J�%�'Z��
��m��a�p(��"l��}�M�B�m�����r����
�y�53ǲPu�
�]��N�a�5 �x/6�a�0"��e�F�����h ����	�iw5�27>V�B�}�`Sv|^��Wz�3�HT�R�D[�Y�o����#�un�ߌ�~�0=r���Hf�b��Q��i��� rjV��=7i��l&��9����n����:���:Ľ����y�\^��
)_7���`�_��~�pS��3��m�	���J���Ya
�<UE�蛆�xy|���w�g5>i8z��E#+���dhc���Ȧ� �Q�\�^��2W�˱A��Mn�Kί�_d��)��*��*s����K~匔!��K�?H��K��7���ͲP�PP>��U�{Φ>>JRk����#/A#.)2�鉮[��*�3t5ٵQ�⥛����/�d蹸�n���#�a�ޘ!ڢ�hX�Ǯ9�q�9�Q#�������WA0�K��ߓ輻qa��eW�� 2-�)���H���3�x���C�P�NX�2a�1��7��=�@�O4G�������];���� Ƈ��{�88�=#[�mm��I)ӎ��׳�EG`�HTA*�����33G��~�Q{�%��j���R$:�57[�}@��嬓c)�\e�g/Q2鮈DCij\����_�yˮ��1�k�Ơ��o,xWs�ir.`|
u�e�R�>�,�L��)��a�{�S��J�z�V�#�2~\}�#���$C�Z�t����l�"�I#�^��P� �_����{+1��s	���������P]BV${:H:t���g�)��Q����o����n�_����zTy&����C�N`�1zR��suw�1�sn�Q��V1��Q�ihU��]���w@�1T<<N�AUer;���N��� �=��vp�r�0����1G���ۨ�f]j�%�'��t1��gsEC��k�:��S��A�v��Y����y�-/�?$��*�'�ѽ����c����?UNCƃ�TeZEF�81[�
�Z�l��QW�rD��_��`z���p��f�7b����ԇ��Mɷ'�9#�@��O��V�f�k����A�Ns�aU�0"������	���ΰ"PD�x��`���B�T���T��L���u����ŀx�o�83��Vx��h��ZVv�¦��ԑ�L�k����XV����E��ғ����{���b�����q3�?˥�<I"]Bx�<����X�p��^>�@��R���K$�����wG���y�7���Ǭ`��v���X�Y)kW�����*c��"�0xJ��������@F�y-��'�d��&4m2#FY���W���Yc>K���Ε������K�n�\�r���VJ���Q;��E�H�ݭ@;�Y"�G�/箮ŉ/��_��f���4~ �
�'s�#8H_v�岡kn�|}\
I
��=���?�*2+��J��z�ޱ�����n�o�ڀ��o�"������Sj?�$���_;��]b��¬���Y�x9�m�Z���P�I����T�� Z����X,�$lD)xy�3>،X�L�1�`���Cv�*�?�2��8��'�|�c�thË�����"f�iƄ��ԗ:�8�0�9��K�(�!y���?P��K%�dTx�.P(���J�9�3��_E��#!1�^��q���ܕ���վey*�]s�a��O�u�\`�Pּ���6M�h����̔o)Nm��u� W��C�������C�i��#.���+p��$�d�e��{��[�p�8��C�o�yu����Nk��C�ӟ�:��Ë>�ǋ���]oP�`,���l��"B(?��bu�G�G���Q�A4P_��x%�P��i���\M)�����ߟ:8A�|1D����^ds��r�pӲ���HӍw;����5��0�t�@^�4E�, �&&O�9����œ��8n�A�.�C��R�(�R�� A�w��~{����]l_��&X䎮��1,@���m�K����
��]����`LQ��oz���� � �D��w#7&��)�8�Uh�{���{ȇ�m�����l34�	p&� �I[O#�:z�7�D���{�\|s��N�r#Z�����4���J��:�e�!��e+��Ϋ��n����1bT���. �g5S�
��3��D�餛�O��� �hh'k��x�0���<�<�D�EP���x���R�-:�H�%m阝�/�k�	?��y��D�A(�o��}R�F/�|�bm���R_��RgO�|����C�ǔ�0� �9�<�ZV}@nC�d������ڞ��1d�����6�(�AXQS8�>��݅9� ���6�}a�u��{��0��z��������d�q�P���X�Ha�S'Z�|�U:�un ��۾= kK��^;�^�:ȗ��j��/3�ݯ�t_�wn��YJ�UB�߽��P5_Ww���p��u����߶�|^�1#gx�HSq���Gk�O݈xNYGC�	V]�mU��ވ�p����Q-E,� ��Uߖ��o씵����)F��/1�7 -S�ٔ#q�E�������.U���3�Jh�#��g����'����(�B�(�S@��a�ɩ~ �LZ�h�����\9�����L�JPUM]� S͞�nB��Ѧ��M;��mbC.�,�vM����W��-Ŀ���@�ʘA.&ǂ���~.�����5
��:��`<k�@l�&�X�k�@&��M��S!�j���S5ש�u�P!�NP�7\H8ϢΞa
�L�����Z��}�h����L�c=�ދ���FB�� &�v����`;T��<���m��ơ��fB����WI0�W������҃�{�})KʒѪ��,�q��nT���Ra��ܕ�-��z�ʮ�7Nq�����T޺o��&򵀕 �1'`O��'U��*�7QG��O���᮳�(��h���gp<@�5o,L9�c?{@~\��S���~b�JX�A��E#��-V��@z�Ci�r4-o�>4;H6�F� �EiI��@���I��w$��u��,�Ɏ7Pڂ�=������9쿼�6LĻ�fw��zЁɮ�%-���?+��>��U� ��ν��"�8��v +�B4Y��X2�)���N�d���'d<߮��Z�B93���`��:�g��)��qq�V�'yt�/�E��Vt�T�&+�$��a�-k���ZPݠz|�"^k�Q���]rLb�^����h�� �y����Q���`�����p���!����5NjߎE�pj��أ���Xm�O�8R-Ĉ���a�Z�d�_"�)X��]q$;��
 �W?��^�����f�M�(A@�u��	�Wa2� ���ͿPI.��͒��+��%��4�]V���>A���DR<�.No簜�O��������!e>bGe>p^�j���#�J���@E��6���ZBlf���7���rhzAb�S��@�;2 �ԫB�y���Jzq��?��t�A�����J�����WF؇-�~UT���l�����R�t��O����i��MiF�JU�Q����dr_)kP�9u@E�ީ>���-����e�U���{Ź[�1_�L�Z��g�)�T���#W�W�Em�����h:����Z����W�4��4�ܪ;�q�Ɗ�R�&�t��;�L�W�[=�#��`���)��p�����(ҳ�F�����?e���](:g~���b�8r�8�y�[���!m�<��t�<l�x#.�����Q�ճ<2�MH4����&��M.{FR�+V�J�E���5f�7��x\h�b�m�ޣ��T$
����gӥɶ�A�Q�����PL0�.,��t�K�N;Z�����׎����:��'�����z��9�����@�Ժ�^�d��
���+��'���U��L��������d�or��*5�K� �&���o���:�l��2�#��3� mEMd �0A�8<D�
V��hl���z�%r�{�>#���ol�C��YX�>|��=����O�^�X�m�G�P|=�/Y+�m3`��H�$�/UXU�t/{� ����Ȗ��#f���sXq1^aM��z"S.�T�Xd�NO�9�^ʕ�3^7�0�!^��h������3"=o��@����W�vހk$�g벎��b��/[�L��V:��UL�qj��w},��,�6��:7��H�ؘ[���!髵(_M{{�g��q!��֞�M�a���}���h���x�kQ�z���Wn��F^=�j8�`�V����[?-%Z��(���4^�uK�M�����z;:�9t�-�kє�Ro+��'�(�Y:�	6� ������aؒ���A>*8�0�,�ϰ#��W��Xf Ӈ]�)b����zh�"epǒ{���N��2�h�t��l�e���b�_��5�>������y�#�p�k~Y���-͆�ʨ �"b�@���дs�S�ap��?9��*��q� �*�����Z��>	��S¿��A�>[�؞�����s���l�BLi��)`��&��.�~��XH�-�'�.����`�ST��������ٶ����A7K6fݲ"%��G_S[�B�,�����2͢����l�?=���v���1ĖP�&3i<��YO�ZG�\r���u��s.i��8���L��}��4���W�E�oğ��e�paKNr'XD�wLH�]�����S�� ��6�G�����e�M`�w�<����$#>�1�hBN
9�?�m�X2�Rd:����e�VN��,�'�I�?�WeHO�;ڜh�X��+��ݘ�)�Y��h/�����x1��u�D:�JO�{{�|�M�߈W�Y�аZ�?��
��(��~ ?�d�xn��A���ժbD���ǲ�7ݩ��WϱUL�Z��F��E��=:H�L���5�)�s�Y�LMyW��~����rw�zV��B����yB ���2??>��B|��b��'��J+\���/9�<0��BT�?��Ϭa5K��E��u�`q������#�2���	�n��6������G���@`/׊'r)y�T���������y���wo?mӨ�eT�?�"U�>���Z˱#4F�[�#�	�L+�)�'Z�Z����ӟ� ��t|��Τ��u_�,��۹ ��Ċ�z�}y�K����a�A�$�˰jX��u�(C��v�(� ���V�`Hn�SQ�"���W^�J�\H��hYgŀ�P#�[��R;s`��B�?�}af��|��M����Y=7�z��6�ry����F)�4�;���_�4	j��ڲ������-�ѯ(?�U	���˻Y�b]ã?���Tz}�YU��bhGY�	W����Kg�U�.jڛ����R|�\
�<������:�������U%-���:���Y!��� 2�b�No�ś���Ӕ�\��A �<)�'� #��芲k��ko炖)�W�/{ج�����QϦ$�!?�z;D��[d�Q����$�y��~��2.�&��7=��¾����:�E��Q�����@���O��Q>Tg��f���-9�?\�(�o�����v-D���OْU�U�IA|1]L)�ygC���h��>a�ufD)��*�s���:�:]3�.��T%r Q��n�0*���(��F:�4+xO��:��Eد��s��.(� J��9�����(:��/��s�C��Ls/1O4<�xi�.��,�˓_ȍ���Jmi<���}˒�F^ä��-�.�h~�I4e�4�I�v�<���?��О����U���;l�LK��h����Ls�;��WR�2����A���"��͊��e*ƒQa�o���U���˂�{J��G�uQ`-B�\]���Z�Æڷ��֥�x�7��!����Κ������:J�̳UU�QM,e��K�e�~��k�x�\���8�`(;��Y����Gm���w�(hYGd��>m^�Xmd ��Sdу�����_t���׌doڤRʬ��-��x�ZP?L!�����[���;�o��h��+��k/|a�q�?�H�H�y�R5�gsW��t��J������&ϝ��v{��X����Ր�\0�~yM�`�~��mJ
2nqb�sTms�9\�^}?yE?5��߬��L�)*_-V��I�����aR��R��l+w�W���Mg�nr�0C���VKF���@����ӗ*��_�<�D�7rCA������b�[�Z*���Cu���)T�����"�R[�9�L�P�S�źde��Ȟ��E�K�Z�9y�q=/���{����<��v�9ܦ�עXh���2I��Z_�3W!�_������Z��*�D�>u���|���-<9Q�������L]�ŧXM�:��;~�j�m�=��Ţs�Y���8�$æ۫"+s/���{B��iY����wƮ%��y�Q��O���b�Ͼ��E:Ë.5�iwצ]N�i�[f�Q7	~��R���K�ށ�v�0��&(Q�e�k�@/��*
?�|��H,2�;mCXL�zxDiuFo�?��e� ����F�V�[��ٞ���{���M�d�kϔh�	��m��-,t��c�W$Ya�9-=`bi9Z��'}(�ě�n%	������6�~klΦѩ[��Vt�M�b��� S�x��j���Rm�cC�7����o�c�H�(K� Z&|eԿ1`��l�S�mYטd7�C�1xcO�vֵ�|���rY*��&���̮-�)X�.Z�rf�X }�H)�%2�2��&x�#���^?�Rc��Њٮ�}�c�D�'`+p�����92�e�\Q����O��u�tAg���D��F+G�D�M[�Ǵ��*by�`��cߎ��%��kI7�g�H�P�x�V�h/J���i��V��B�&�yvwK�X�~W,K1�	4��?T�)?�/����KC�JG���V�c{�����l�H�x�V�C2���ݯ;���O@�C�Wc}����Wv��]�n�"�8��g�jؠ3�0�uǱ�[�h�w����2���;��9v�L0&��A޻aH��ih�°}'Y"
�쁇�2c�=7{|���z!��C�(�E��J��2b�)����bM3ء�u_Q%��,.;p��63D_�J��e��/x|Y�E�����M/��xn���:oRZ0���
��Ej:*�����y��Z?#,J�d����"`X*��&�n\_&�O�S�Γ�L���9a1����ka���=#�;I����&׻���X#�"Ģ�V_�Jcӝ)+;o3�bմ��v�l�jw@�G��rf�#��;+G�wm*�����wD�Lg��ɝ�V�`��w�ߑ���g��,�ڳ!TxzQP9�XU��.��F�l���6�^�qf([��[��R6D�,/����B*o513�kv�����kDr�s.x�_r��!�ś>��͌�pM"T �����^��x��Kb#�ϻ]!�ՎA���!uL6u�ym)���:"ed;�cPe�[=�G�����B��8B ����-P|�%���CF��_4��K�X�VId����7���"g"��������kV�cGང�\X>Q,�c�Q�=����~�i�_I)��W �ƚ��OqPp4���!C��i��@�<��`8��C�~�d<��:�r3���xٹs'�����G�O���2�t��W�V�GA�+�M�j�*`��3�7L�QW�/��'�2����L�=m|:�9m���(E����j"�0906�)�"�U�|rɐ�Z6;w��L����q8�֠�-�M���?�/Un������sh ؃� |���7^AԪ�b,�`�BX�ĚR�����oDV!��Ś����\lď�% ��m=l���fEU�ǫ��3�5�����AR�����"��0���rmR*�t#_�%�R��9�Fy����D��Z���Vĕ��0a������u�Iщ��D����.���Jl�~˳��"	.CvShì�[������_��v�73������Ge��NOm��Au�[W�?�����@�!jw���+R'�&��+�@#M�Q�єm{Y�*���АlD�-��n�U�D�MC�Q2�0�N�Xӻ�OQ#չ�U196�*[���8Β�߰��}������m�L�H���7kudg��L^�Dh�i�Z&2���H�b�9�L����Y�b�Z���I:F�}�;�}# Jzo!�DQ����&��U�N;�u��:�a{�w��k���I�p�|˲�|fq��D�����_֩&����U5ҷ:D����  6*R�����!k�_��Z	�%_=�9�U�����vfc�2d�V���5c��E��=�EZ�TƘ�w��e�Ê�5e�Z��A'�j@������h�&�=�uI����9�ũ�Y r�����1��~�vr2��L;��h�;��m�~��TQ�)�7 -����E�ĉ���	��/�X����KyǍ�U�^d�V�����%ۣ��b�G:����v��Q�C7��]|ɲ�g&�.P�O�ߦm�F�\�q��#���<��	gb�$��mEa�3�l7*�|�O�'#XK_mO�����ы�n��1^�6�Sӂ�]��m
%��o��`G�*�C��k¹G�*�?l��5<NY֡�����k��X$D���R��-Z˲�h'V�&�Һ���������GrU�}y���Rӆ��HH�ú���r�sx��! EVu�x�2�~���1�b�0��啦�K�Sp�'fyn�u�uS5��OB��k;CV��>i����͠ˑN_�".���(QV�c��� ��t`1�V� ��8��%��B[�d�3uܪơ\�EV�����π=)#L�cR(G�����e<��6�w�ȒE.6�� `7�9�N'�E�A�<�<A�sB�F���o���Ϙ�K
����7�2�OTŬ��A̐��-xaK�Ri�VO[j����E��;n��؅:��@fҴ'�Pr�"?R���~U;��2��c�D��_��Q�)���E�̂�� M@u_�J����^y426JM ��7��#��t0�kbS!�m��G�������P��r���[���蛽�ᱟg����Խ�B����p���s�5y���3�j~KJ1+>�%99H�����yv�y�f�����)YE��`��v5HY�.�S)�y<�BҶ<A�4����Ӝ~1 ����B3�Z��q�����"m��{�0<`$���\��O�b��W6S�l���X�h8
���!!�b�W�2�Mqጸ?Z}O?�¹w�]3��F/��	��&��C��@i�����Ҹ�`�<�p��w����]�8|�AĞ�%�`�=!A�u��WV�|����5%�އ�ek~\��9��7g���Z�x#<"̃��1��F��Y�k�f����xr����Z����o��\�[Vac���?���%é�QK�5ۢ;3o{;[c��sc�/L��L�����n�4�C���]<�Y�D"V��ӧޘ.���;�%�%$H�ހћNmJF��f�,�C���)f�w��c�`�¼�iz3K�/'������y+��a��� ���LMJ·�.�?�8w�)z+�;��V�Hԏ�>�����J��F@\�����T�}�ǭ�P���@��l�`PBPr(��A 4n����I�>����Ya�G�#D{ �c�Op����G8Z�=xP� t�E�g[�T�y*��{X���U8���[���f�+�am��P��O�Bg��}�À|��9�z��"��g�`=)I�[ҏt�P�c�zD?dB���G|5�+4�+/q2xU��N쟅��Q�0-���� zc�i�&�nj�S�[GV�MӢ��4� ��'�:�SX���P����r�Q�Jk: 猕7�[��a�Et����l���7�k7g1&�=2�YAK�I3��>L� �n���ےp��'�tZ�7ux�ij�}�2�H���+۬�ԍ2�����/t.DREJ��*�"jYd7'�ڨ@:�_�io���1@\�Q��AW�Fa��yq���Xz[d񔰢��G�iJe�J����=��±��I��fn��O8ǆ���m�mD1D����0��
^��BO�c�5��o;C�$G�I=3neNrc�+MM�8���!�c�n�qS��7aޚ���*�M�Q���+ �pT�v���쫍�K^��g�H&����,F,�Y\=���R7>�6O����K)��D��qfG���R1��� ���8R�����1��% ��zF��3wU��LH__	���[3z7hCKV�Ʒ��[-ծ��	���X6�:���+�FW>���ѫe�~+N�H�5.��'N�3�t'{l]-��_4�Tȃ� s���Pu��JU�*ӐNJ�ւ~��m�e�26U��Y�x�X����,�Y1��|�Wgc���5�(�G-�V�pY\��U`�a�j��
G�C�b�L����O`C���}�aw��	�.�<4���oa�d�ݰ+�el�tW}������^>��=�Z�F�ͫ���wYVL��JO������z����D��Gm��_X��/P���°=���e	�̽�$��'��#jea���O���C�}C_aX(q�Y���&K�4XwoC����>.m���f���#�x����[ar���V�:�̑	Ő�A�	��f����Fxu�O^���~q�^Z�>���N�?;q�/�sV2�ݸ��s��45ލˉ�@b��3�[��<nqIʧ��9V��9�����/�(���Ig�.����*}w�+կ25�lFQL�����F��$���ER�4�H�g�*t� �m��0�F�A�}}��6�T"��-���Eq��1�1!��K:��[S�7ڴw*�4`sh�|�E�f[��E��Cޅ�M7�z�C�UB��p���o}͎��
@�����w���=�� {�HA�u����ȁX�!���_����vw�ţm�})&��*P��&���4l�����H�^��V^�38:���ZT U�9i��l���p�& ��x��]Ϫ� bW�����C(Ĕ.����*����Ĉ7��T_9:��%��U{�|7�p���0x�
	7ގ_f �>�y��|�D�t/����m��b���\�4]��[���̘@��$*Rh{�ϐ�3��m
W��}"k ����8�B�؅l�?X{�!7��k_pۍ̔�s��HR�6�ѭ9��{_(����INaB����Q�^�#h�(\�n��hY��Q=��V�D�f���.��d�r3&���:z�(�մ�y���&)�3_�-�I�b�����;�{�@ �?��=T@Vw�*�{���*2Yt�0)��gH�x�5���ѮD��\�ų�����.e���K���(d!>�>���B^��4VP�p�� ����zj��<�gҔXL��e�z7w����J*���[�M%�R���a�η���{B �:q�\t|U
�^��Ԁ���]gd�Mp�y���������~��c8���|8��1 �������W�g�pr�m���	 �����[c������(�7�����)�(�BZW˫~:�'S#���	�5%O���'l�g]#"3N`zX����Z(Mx�r�EV�6X4�1L��ɬ�"C� Q�Md�g3 �(^ԣM�>v�z�"�KihF�"!�0)It�> )�xGF�h��Ot��11"�3m��-xN��T[�Ϸ���߄'�u���o׬�ZHz���h�+�/�����P�# Z>Ѷ�n�\���It�?|�md���y��/?��@�\V=�~خqh��������Р�5����]���?��54J��l��ik�V��F'+y��-�3'��am�_����V����E�u��dzf�'&���U�M��zv�����~R��o�H����2��"(L�>Ǘ��>�A�0�
jJN��v�aG)eV�k�`�kZ�������|�=����YF��.�S�EY\R�UD���r�8O�.JE��ǬU���i$�v{i���C���^����B�h�s��T8�@��℅{S�~l
�P<��	��<شF�φ!�.ܚ5
<�Pi�ڗ-L�H��)�����cJ%1�w��E@���$�c-���f�"[d�碔`������zQ]��x[������c�cH��1oo�3lW����@a-�pw[����
��hYkgɥ!J�=a��<�������IVX�d#(�pň Zo�ZoJ�с�0�b&����Ԙ�܎�iD�fCC6����U^��G�Ax����s0�����Cp��+��W���?,�G�ۈ����r)��{�!���P9����΂�����|��U&Q�6$�D���v�'�s��H�Y����;���^TM����k.'`k}wi-ܐ3��������$j4�U����Mt�+[Cy�����NJ���˖��m85`H*�J�Q|�|V�pPB����Y'�x#�k>��f����]���E�`�������s!��P�*('H�$�N�
-y �7n��1�j�jN�z�7 ��I����.2u�~�vqi؂g�2��m�'�
i�4��t��M���>�7�b~�l@P��~XJe*��:��,d&��5f�����x���V�b*Z�	��N�X��q��
̍��-$�6����#&��G�츲v��+�n`#�k���x�ɢ���.U�+Wi�>n�_w��c[PKl�4�M��?���4�z�e��<�.�ʕU���Q&S�O����xU�+��؛�/]���إ1�j��(<�8Z����Gd����X��$]SL��|]_���~ǹK�>{ݿ�����d�������5U�|��E��<!�B�-�Q'���U��W�>��c��0s����a�G��	i��xҵ)�k� Y�Z�H���R�
��$�^�}�����IWm$a����?�B�\@��JC)G0��z����Ql�.����h�����)�?�A�3#Hp�PH]���w	p���zxmxR��?�/H�ܬ"���<o�tN�iL����\��"�!�	m`�<���~k�~+���{�J@�G��}.S���u���d�&�31�Mg�kJsh���Z�����s>~��ܑ��\�Z�:7`�Kz��M�睽?��vjo�PQb��gΫo��J%R#]�V���W�3y��'��5m�Ȩ��(�k��"���4�� nF��Ee�j�TD��
S�p|9����x���Y5�J Q�n�'gP�u}R�l˃�����ԘI6!1���U��I�LD(�X�c��JXC?`���Odt29��f&�v�N�|���.���^_�������kD�rn*TV�m&S��õw&�C���I����cɐ���i̍�vr\�*~�Խ�;����DL8�sǧ���7�s��t��_�PfU-rW-0���ɾ�/W��С!��y�n���Xb�E�J�R,�,�{���0���MR��K2�8:~�� �R�S�=y�'���wێ&e��0�-�.�0$F�.��2E|�d���[:�B�FkN�S��-�?���³���κ��{������QsJ6lEPQ�b.���,h���0*�W�Cd�;��i�kJf	�XJ�MX�-ݿO`K��!�hf��k@���:� �8��~�o�!���<�D�ꦍ�>�1F�o����x~�
蚱��ڑYIl<~�'\��'N��<l�]��� �atH������) �@�F+aO�]/�h����Ӷ��A�g��Ӕ
(��$3�;���ԟf�r_[N)��W�J�+V�]��{K���K��{8��Za��g,mV�N;GZ"h>�5� ! ;çeo���»�=6#<Ob����+T���U���sf��ᙛ<D�T��qcãY Q6΢�D�J �E>E��Aml���c��� ��fvPV��2	�Yǒ}R%qVo�z�q`��D�,r��TUd��)hG}7(+���ɐJ�et(P�����|�5?�����J~��?�oAE��L���qOp�`d�7�:�u�ފ��E�'�!y7��3$縆�G�����ʻ8=�v��=�/1(�;q�%u��;)���]lԶ�2�t������²���ǁ7�a��qD~�	�Hs� M>���Iז�B��#W����oT��ǚS���^�V1�ᅠ|��F�^���$u�5$��dm�4f\nb�� ^�X�����n��
���A��S�����܂��ʟ����R�YKpl	&�f|G�a�+Yd�l�j�
�A�4/�������ŜOs�[Ԑ$�(-�O&Kb�g��)��z>~A��O�>��7�F�Oo�����_� Y:�WNh3Rݥ>S�䄖!�yd��ˋ���Ĵ���}���%��%�._k5�i�<,��8�Eo����91�vcӰ߉�Z[�oc��l�O���1Bc!�CG���?�7�� 3�ʲ�(A�
;��E��O��T�*ѝ�Zvً�>�})��L��(0*>�Κak�%ӷ�m�7�/�C�fJ����P�\%)|W�}�:�&����0����d��v1B]��T[��aJ.��Q�>�p�Ӏ�LKB�f
oD��|*4sQҭcƁ�� �Hd��v�qD����k��EZ��+��I�y�Ra���c& q!|)C��f������I����7�Gn'6�l���Д!���Q��N�;#e����d���*&�SDO?t�z~KY]I�I��9l�f��"�b����ɷx�,'�p�h����u�{rV����ɥv��X	�:Bd)tnu��uO�?�������ƲP�J&'�Ee�H��R��L��@�}��ܰYfIh�'=�-f#q@��yf���z���]��n�Z4B�2d���塠��k%&��#��L�ȋ/���d��ۀ�N�<��6|L}0
�|�I����_� ���t+t�K&0}Is�·�^�!O(�äou���0����'K�^%$��Ǳ&}ǂں�oxi�|q�P\��9�F����{HȆ|z�|��OK?�Z8�8��㉰]�Q�}3#b?���<L��͘�1�@tWMp����/S����o,az��s�*ڹNJ����ē�c��R@��hM4���דW��Ļu�\l=&�� mK#��t�eD��*f�v��^��ػX'9�Ɠ[E�a}^7"��]>F�����x����8�rIs��sx7#GCv�f-��Tv'
M5��ʚ~��nR�X��4�M��u\~�Ua��x[�_g�8+ lXş�^(J{�_U�s����W1n�8|4�g."���Xb�H�[0"}ճt+��^=.�� ���̅4m	\&d�P{c"���#�_�J@�0�L��<�Lc)~�s����7��];s�����
�r�f١�w����_03���Ƒ���e�(��"$��oQk���ˑ���D}�#7ɗ��υ���*O���k<��M�?D 1��F�֋>���E�Y�zk�%"E\b�-�S�̃��:�3�vu�ͥ����rT��Y]�/h�*��k���'[�]k\�c��i�䒓&ղ��+ �����?P::��0g�P�~ߙ�^6��\&�:%�y��N��"rO��1��C�Nn�I?�� S���8��j-�2�.9*�kb��i?l����^��Ɍ�oE_�4�ƲI�d����0�L_N�Fp���_jhq'���=y�tN.���&��F�)��ŋ��D��1�Hk� ++�U�P��+t�6�?A�P)�B����:�Y`z�7D�"@�2���̕��囤ţ��Xv� ���w�ji�u�F�Z��߼�	p��#l�"�g��<c�)s�n�2$M帎�:�j�iӜ���	s�]\ӵM�;���Y�|�4�s��:��)� ���1S<H�QԚ�AUh���۬u�ZcWE��J~ۓt�A4T�	~����`;7�8u��3-����f���w��>������W]P/�e:[����:�2��l*�7����;:r+3�`~8��:{��E�T�Dk��j^4Ni�: ��3�b��|��囐*�
���ZL��q�])'����W%0l!l��=�!5����yj�8�p����%��iW*�#� x3��G~	��I[�ݯ��?� pQ0#,*nzZ�J|I���0�*4�,��^?�6�ZO��]��-pT�#i�}7ս��ۍ/�S8�ڊ���I!U�$p��k{�����Az���|9
�qj�$>2�������Q֔�j>�^�1Lɯ;�l�P_
6�����⼒�����&�ٕ�S=����+�����p]2j(�<{�������gַ�>!,��K۵�
{E�_d")d�_���������$;�N~�Mx���=��79PZL���ƶE�v��4e��3@	8��63���4
Rcc`]�&�u�p�G�G;�C$��A_U�u�}<�s+�;�L"�㰵sd��雃�z~�'w:f����6��8� �J~#�t٭�\�Y���b[�Mc��Tu�-&0� Q1���J�y��rY�0M���-�/U9܌� �dl2�Iڸ�Ą�z)����a�ax�?6�9 YU �Ž�Y\��\D�WW�lB�&O-�}�X@WNN0��������%w�\&�G�XuY�La�� f�Յ�NՈل(3�l)�:���3v�V�~���g�zW��=-����[��S��hd�o�*��+:���|����-ۋ�M6.缃:\���R�9��ðe.+��~|](F*<��1�aWn�)�����q�fd��vQp�/wGk.��n�n�1��E��G�����aO�?s�L��gX �!�d!��gĮ��5� �H���L' D?N�DҢ���
݋��n�p��ד�S�Ŝ-�n�گ�!|��;U���sv?���ei]�F4|=�Ն�81 i�x�(�l��ƍ�a,4!%\�F`swe]I��
����z�&˓h��ft{�K��u�[4J]�gzS��2�b�k����r}��l�n�M.9�3k`�BƎ����I�������i��b��.�oV֌@��(���aZ�X��5+���An*�L��p-¯�tq��^t	��G��^ǂNtu�b��;غN��)"HB��L���F��8>h��9�"�㣡�>�e�P�u��$�����@RW�ڌ@�t���܄��D��'��c^r�g���尔�%�zT�/-ǻ� �h�� �$�0�+�BC�G��$&B�^y.Y���;>6�~A������\e�E�i>�R������bF4q��J���D5qO^�'�#����D� ����~�P�1�X\�,�Vޗ&�|�<���z��,㾰Gy����6�����5qC���A���i��s�S�*�0yn8LZ+��'5-H�\(0��ބ"����$k���9�<��N\�aϭʊ��M(l��k����~!��VR�P1��M�H��gAD�l���Sߒ����dt>�5P�1����ی�6������ߢxS�.A��щ���zq]V)c���}GE����㣉)�
X�Q��{��Swnzt'Od�U}[���ǳ���"td�k8Zd$�3\�_Ժ��[|Z^��(i�l`�[cs<(�;��/�0�5,�H�G��ey@��b�����q�2܆R$� �ݬ�^��ۓ>��FNGIɠ'��^Қ��#/.ۺ@x�G
D�;0e�^�W@��l2韄�|ʌ�n,�kl K/��E�$Ȃ@����r��Md$�W��a�~
�N��nJ���վ���<B2��B~J��B��9{�����q������7��ܪ$2%�m�K����x�����(��+c���?ƺr2*�3aL��^�F��~	��a)�t���I�g ��}���x��� �('��L��-9Q
xO̓[���󆮚;|���� "�)���IQ�ǧ���	�v���6Py��2�j��-H��3�ۜ*��0��*���� ��׃��e��{Rs4��\Dy�
l/h�Dը�է8�(\d�$O� a&I�"Q&`.����Qa��*E���40_O� ������~~:�;��@�F�-���/>C��n�I�e�D]%LMX+������8�Bb���9�GV�]`ŧ��%I�'@�]Tc�l�}/��pM57T�!K�v���/ug0�������V��w��s��>�j�<�$6�]�7;x���,���ֺt$���#��i%$M:��'���*�f�bE�f��=�ZK鎓]dZ�X^S[z�kS�V�D4
B6���s��w��������U��2	�b^?0�������ʘ���L�ҕ�>����5Q�M� �i��D�w�s�,��Wy�H�鸖;eJU�f4B0�*��zّ��Aa���:\#�NKi���4�)�ޣW=��F(�79�?�hZT�ᾛ�R�W��Y��,D��h�-��گ~������W�O�g����,�[t+k:�a�p&IX;��;��!�"Ai+��wt4&LI!��w����˒�p�`����%'�^Njx~b�@d3w�]�6B����-�7�eF"ҋ۪��(�g���4�bqhIA-�A�T���@3�RpX�"�]:�
�:��y��&���R�ʕ?�dA?�G��j�D�b��?���a��[�%��-X�$�I�6�"+��A��8:RI����v�5��Z���9��J^>���JD!콄o�C�质�7�3n[���8��y!�n9�d�����lm	bW�C@Y�(:����Hn^�E}������*^���&�'��`���^m�G�ҫ���;D�CU�!�$�m�+��PG~8�>�DI-U��a�*%)�zr��~����z¿����t�)���Uw�oTɹy�}0ʨ�����'R^"}�U����I�k3��Կ$
�lO!��m�I��&�e5�0q<��N��8�y��<@u���.P�+&ҟzN2p^���q����AO$�4�fo2��!�ǈ�W�s�	�X~���s��5w���I�����|�Ȓ�*>rU�U�Mck'�h �m.0+�I�w�	-�c���2��k����A(��m�*!`CY�ZM�"oG@���[��%fP0IM�y�|fF�R�0gS�(��ڛ��k��K)1���G3t����{�����{��Ep&�I"b_���_���~����|���Z/C�`���,���-q15�7BR��}%@� ?��ZU���W稰N�Y�[Hl��ժ��;?�2�?2;���Ιw6��^yJs�7|΀��ڥŶ�W��с��왑GgW3��;����8B����	��#� hF�ad�wN�3�p��Ҵ�!��.W��QV�ǯ@�c--�T�M��_�	��	?��<h��'�k�1���{5��v��Mo��I��&a.����=�����0�E���������H,r�����ˍ�é�v��(�6~��)<��íԄ�ܘ3r)�p�O�rRNP�e�w�)aXx/�B�-o3sn;K�G���S�P�ؠ�e'3�Up�PtL��A؆I{<�[s���1EN��!)���#$F��o�ie|��v�L��]�X���T��(�z�L���oo�D�\:D�G��3�����d� �h��JO#�p��n��zc�Ru�o��:u��W���V:�"e�������V���V�V�X�Βٔ�lQ�8�%���;Л ]�` ������ԫ� 5����P%~;�Ӥ ��,���y}/&�<�͙2 �A��i�AN�J�5�9�&��3�G�
��hZ�����F�f�ʢ�؂�{�7���0ik���蠝g�U�	)�c����{��W���*u�Ɩ�f��)6��Y���YUQ
\?M�:��d7�}Q�g�Q/�%
W��y��K�'���_E ����Ӻ�H�P)�F�ك8��%��,��#p���Ϲ��(�}�+�7m��s��|ᒟ�yi��4	c�ߖ��u.�n�/>r)e�i�}�w��h����ꖔ(K����a<�4{o�?�IM������A�e*<�(�ENY%�nH�!�TFɟNU/��?h�5C,c��5�فL��*ȿw�u+��N?��-0��z�c(w���su���T(U4P�
�1C�u�+d�I-�Nռt��S��0@��!��j&
�+㠿�/�f9�;H��U�����a�&����𚈶�1�)t��kdZ��#uapnDY��#��r�?)8R)���Zј޺�2!�"���!�Idō��� ^��$�����35u�8��y�a �*����-�l���^���!;><��5���k���URM�Ũ�G8D�k�%7�`�GC�c��T\_��c_�N�5*s_O7�PK�h�#Jo���S����X�r�~�%�Js�KRm�ڞ�����ʧ�X�)��@Ơ��]Ta�i���mϊ"��*#x��aU�Ph��a�`�0�;"(ag29�l�V�f���U�9���>�U��M��=�쨥p}ڂ���i�����b��Q-�;k��p��� :Pj��� г]`T�q��)�5�Ri�J����7L�l��{��¤ĸ�KC�}�O��8�M�Ά�~3�a�����YC|5��x�Q�
�NO3�uW��:+_C���2$��e?�zݝ�������R�9���4���|'�|;ѥ���)�o	])0���Az�/ت%�'U%�Q�א����9��&
���	�O��at��ң!NӼŞz�o�ՙڸD<�C/2�y�#K pCvej9�^��>��`i��v�B��a��W�."z�I���p��F���x��A��#�
ZTWe9�ܖ�zpx��$H���zm� we�Qm�:Z�n��%l7~����Hɘ��e��O�]L�����V�\���+���ʗ1���������>�,�Em����y�T�k ���vꋲ�	�XAFՖ\M] Ln�"�%>��'��I�/��i���aCC�:%���h$��U.y<i �ʬQ�qA��'�)5�������%9��>jh-G�;��`��󦛒��9�5<K�EV+O��?I]��F+��ǽ)+��+���+|��{��[X��'���J�d����h���r�)�stđ�Z��ä�.gd�S[iͶ�x�4�Հ����i<��kB{��GVՅ�{�O��+흉Mڪn�?�DuT�z16��L��V�y����f��?	���jQ�xĵ�xX���G���'#���B&/$���1��ꭔ���� ��l�JO�IL� ɽ��(�ӌ������m4?��pF~���@t9~9kS%�sa1�~W���Z�j��Hb1qo{��*ΤM�Fc�[�2Ctצ�[���ˬ�)�ZK��y𼶞�rQ坲k᠐�)}]��m�}�1��l͎�|c[L�,]!}�&s���4��Y�0��hc�2�����^��@X\s���1]��q6E.��N���F~�27���"����\R+%J�rj��-�\O��/ j3�c��7�:+(��/�ڈ�M�=�|�{�>p�葲�|�9���֢ݑ�Ub��|I�+������a���c����)5�n��e�{�-=綹����f��r��^>)����/l]�-)2�8)ͻ2TT��	��#�� ���;��~E��9� �ņ~��[� YW�,:+���<U�?kG�6����S|"y]�P�7>�)��k��kU�_Ű��if�N�������n�܌I:��j8�5$TV
���n��[O,a��k��Ɵ(�2��-'��>�ke���9c��<�[�>����R��-�J�-M^b�Du�幦��@5�9ߦ*��<������<���jZ�lvx�á�d@��Q ٴ����_e����~\u�m��!Q!6v��:���/��O�:GUYEĳ�gm��~V��8Z¢�]r['}�G��t�=���+xQ"��ёH0�]�&Ԝ�+V$��*pU�N�2��a+���Ó15���Uo�0eVak�[��ʻ��Ms�5ݞ�@GG����P�"Ӗ]��Ƅ\{�h(EX6��v���V�A��1��Ͱ�i�(-�~d�u�__%�,�T�$�)q'����ռ�9a9���e�b��	I�â�]HO���J)z>�_�	��1����+̔��0V�c5����Y�S�hF^��+�;
k�DTHyh7��b�6TAr7W�BN!���_иI��y����߲װ'��V�5�!�8U3�+����n�>������Q�C�QC�,k��`�#c�啖�Hb���I�p�N�OyE:~?QѨ��T�5�����xB*�}n*�����a+�6ʗ~���]��W=� �6�"�@8k���������?�獬�8�9��1��n�G��I�<����)��U�,���ja#p"H�R����N`'l���-HD��Rт_'i۷���<2F�LW��)�%&m.nf� �g��Y&��5ܳ��ib���JI<�5���S	��+f�Ivg�pD�ں�C
�D���]�|yo�T�NzF��}�F�H�Mޝ���"�{Q�o��N�~v�E2�TJ�[�raBP�
�h���!��ͺp�,5��Jv4#�@���V�O�2;�G��Sn$|�4�Mo;:����m�,�i�k\c��i�K��9~��;88l@���C_�^JT�Q�ư-&�6�f�>���߉�.{��hw��|s�2(�cM��A��ϋv@n�a�Is߃� ��c��Z�a��Ͱk���|,Q�V==���hI�άR��͆䳧�k�x�e���hOJ^��Eڅ�uqg�-=� &������k$����3#T!$�x��j�3�ൿ	\�I:ߵq�%`�z��z�
��`t\�=R��E=uu�OV �u�O"��a�a�Y���1�3�x�՗[S�Y�,�P۸���w��/`�b.56͎�a�z�@�h�K d��L�,�k�x�w����2��ؘ5�2isD�dxNkn�*?���j�2�tܛ��I�l�DT�i�5�̊b�%6L�h|75�6����V�5���~���Y��U�����@��Ab�@�Ƈ�([+챾kt��y��L�?�qe��n��cK����U�+�G���r�E)����s�U��L�W�_��Ȓ٫�"{I�{*-:S�%P��`�ac̙�Y�29�֢��N礍��zE �8]�1I�7��|^��� �I#G����u� � �6��n�����J	��I����Qb�xY�-ȹ"�7")#�E1��Ԅt�������\�����ŜQ�5[�T9À���{����X�n�E����py��St�6`+)�.>qY��:ꏷQ�y[� u'>����G
#�jY4�li����<k��6���]��^�Ϛ6�?�`�C\wz��T�1f 
��8�
��B �虝�A�&�}ȸ���F�Q��J��4yq�Z�A�H�n�;��)�
�Y�rF)�`Ty�Y;�:�x��u��ְ�B3�Cr��sd���]�������EϹ7CK�f��輬õ� s����XN�Z��k]kD3E'�^+;��P���e����@�zv�4�L���:��J)�W��){���8�Hh�}L���&��E
{�/PJ�x��4���8�سh��v�/ҧכ��bg�¤Cm$[M�@��w�B�����BԔ%����\C���?X�[ܤ,-�	n6����4���4���\�%6v�NXg�(�ol_K�x��c"�y���-�Y[V=�vԭsZkHq(�M�m�2�qDߢ�a7J
��m�;�rD���q|��w���w�5a0��A�AJ�(p?X2�הL�%?��=�>5�#ta\����Q��I�����ky٧���f��]�Sqv���/�ąx���j��Ԉ�E��X qX�����H����.�<��%�몧4���W�IF;PǇ��!il%�}YK�H��������-:햽!&�ϻ� V�^T	�}+�Gy�;�{[��J�0��鴤l�'��L�n�1����Ż�:5�/�\(BKI�a��٤�[��7�f��/`�fr��c���x�%	#|�g����?�ihJ���� �	#>1�<�ݲ�m�8��=U��P�dM sV�@Б�Tᦡ!�}m���L�ƢJ��Ϳ��7m�4
l 2��n���+����V8^��ǟ�d8��w�2$����<+Y+¥�ftnz����� �B���~d��'�XzƧ.�a����I���r�f��z�6`�o �ʈBP�>�9�Y�cs�bv�"* �иV#�eHCwꌹ�u�a�ȿ]����MN+ƒ��f^�������A�C�U�KڪP��f�"�zr�!�"�� u�e�#�K5(O%�D^�A�4�v^=$����D"��sS�ӆ��6�u��w�Y��Е�t�W�/G��VFX�;�E�:[w~���#F�v8�1�T�_�]��C�0i������.-�P<�J�K���Ȍ�v�W)����EX� "B>���UOA�CCm?��CG�inn܋�y�,ue����/�x�	Bb>�X�,����xe����$�T���*��td��ǂس�/d)zT������*����CZ��u��O-|��;ܨ}�$��p`P��|�}��C�7U̗g��H!�����#����1��	�cḏ� �m)�A��*@��Y��fdy������r���drt�$�2Aʴ`��S!�&��9�d ��b�Х���n�}o��$RrJ���C�E8)C	6�B�n�h�?Wq�h��������J�:稫�q/u�_SIT ��dʓ{� 0��
6#�L�K��D���5 ��Z�?(�9�h��b�y2d?{� �н��T}���x"bx5u|U51�q����@m���ZJKXV�7-O�J�F1�hIB�F�od���m��"�%��Na�	�H`�=vY��Iq��}�@/�Jjn��5��?�]P�/�u&z/x�NWl�A�,�&��E�w���R�3����$f1�/�C/�,�бX���A��I1}`�j�V'T@9�}I��l�^�^�o4�f��P�(�F��v��z����􌕴3��~b�~Y�O=P����1l�����R���%�z-KZ��Ƈ+��֠-B���k�:�� MI��]�� F�b_`�7m���ȫǹ�=Xf!��pP��䈜Ȝ�BR�$C]d�;��e��[�R�D�7��UWm��H��qd5��uvK$�7�c����ds	���g���P��.C�iE
ћ����so�}��z"��~u��Q(�O���0�\��W�0�p�kpG5Y�2.��h!���@���N ����->�
��&���y �P�Y5��fn[��/&�g�Q��,m��p�*�}��}6X#�?�_ 1�܆���%�	U@2�G�}oa�0�ttwzme�
����WdXM�$vQi��C���1����U�S�fó�`�m��_|�))}�����-�����Le�c�)�m#�xĻ�&���V��l`3g��k��q��>�r�ʛ?E���r�~#Nɓg�~���`lF�>�A�m2?�C4���u�Xm������9ب��_������ԥB���L�dۥ�����U�'���˼y��)��Q~�&���\��"�(��|�В��/_?~iw԰QVV��ω
�7��n�/��C�Io���Ap��APg|��6E\����h�ʔ��u7�|+m� �NPC�q��v��糦�z�sM�Ҵ2��f�p�A�%��o���d�'�����v�Q�'͸Cv%��D����u#���$n��e�ly���|RJ�i,���>eEI(��P��u�2�:q���(ʟ�����5�d�]�P�gs<xN�O@�h����t����
f}���h2���۪� V�vc��u]aW��'�?~8����RO7��)���F��_�����.`�k0ϨXbM= Vq�!��b&,'�k��#���I5�JloA�����^�'�8{�J���_ӱ�@~ɵU�f˭�"C���ұa�6S�S8���aF��G��~�Uu�ƨ3"\�I�Rhg���J�����I�$1hA�����1��&�%~1S暽Ua�7`|����ʻ���,��w&w���5����	�X�w"���/a��tc�ۭI_�e���!����؊��҅R�`���?"U�f��Y>��8�h�M�n�	r2��h-�J�7�����3\�(�=oxX��=#cz�	F�k�8�H�}�$U��5h��:��y�o��ǂ���:��x���k)�R���!�К�$�`�d|$��ڛ]R��[��Q�`�P��i�fy�Xǈ��N�-d�S�J����<�s��U���V��ʄ���j���a���V#g,�����GL�F�:{��4�s��q�b�k�{���_ҧ@*�·_�EF��d�ޕC�,�M���{���.��VYLY���1�,��1�-�;
0����
͉Y�j����Q��m%XY�e�#��)���.؇̧|�֨��9�'�ڪ��+�焳�^�S{�q��y���w��+'�|���@\�0J��f��G`�Y>'�Q0�T�w.S�r�|�3q�fh%ׇ{����D /�������'m�U������=n��k���m瘕J��)9���k�/���H���%CTG�T�z��b�U<�u�Hl7b�Y�.ۘ,Y��� �_?�kҚ����Ij=9�)x�=�lb'�㽆�1�60YF�h=!oA���G����v��7�e�?Ȟh�L��ǟ���^�t���Q�T�؝�9�{f���ˊ{S�Xʟ�s��u>�����7���=�mk����.AT�&�rLy�jhl��C#v�}��g9�q@��5T�l��Vܓ;�S�Y�.7N���u4�ա�?w8�s�l=��0���C"��d\VS�yoz9T-��Ő]���q��Zğ���
xpN����؊^S���t�%�'���tS����a�a��� �b������ly�On�X^�ɦ6W\g�K0I�$)2T�ɲ?�y�������ouL�Cć�_]"���T�Ulz�9�����~���%�Qn{aݦ���7��cƉ�~�%5N�rN��!`j��0t�h�X�^&���G�L8�����a�Κf ȭ'�'��u�
�S�w�r�����qC\(��=�-��l(Ps�j=����ä@��y���|7M�@��S�f��2�b�"n���Ю�+���J��Ź}^��V��}z0S�M���Uw_�V%�+২��)����}��W�B�M�e�Mb�7�_���A��o�����7��x��A~�ښ�	�[Cg�����~(��X-��X{;3346nmU��;`y�i/������]B��iN�H��8�L?Y�w4As]� �491Dgzӑ7�^fS���B�ڱ-�DӖN�h���Y�`�?�S�<u���
Ϥ,��\F������A`��H�MY�-j^Wl�_uz�����ݘAMM�Ҫ���PW�iǦ�F��z�Rd�G���ņv;��|o�_�3p8�?l�]|�w�wr`���[����q �o������Q�r���,��
�몃��.`�l5�~�ČȆȹ���[�(����~���yW8)��v@H�O�B{����9cu�S����wۍ��(�Ø��'@;�u�	4�.��~�'��}2�րt��`I�&�05��� b"�v��#g��,�K2��q?�/�!%�B7t9g���&y�P�� y�֌��=j�A���
yT�4ڰo�F��;����L�E������<4�~�K�����P�����W�
@�S�yN�������	�qN�>`�7"$�'⟽�5�"�g���x��%/FQuk��bה�>���Ͻ��;��b��� �>�h�؅��^��Ш~j8��R'D�c��N����h5`3�/}�ܒ	��e��4P�bHq!�J���������$+�S�+a%�E�E��1 ���ҺO�-Vmo0�m��#М*w�s�Έg`6�ҵ��#������7��\�\�TL��._;�-p�=�xd�p��;ۄ
�`�&�89�ɢ�&�6��
ȣ����{�b�vyT���\�����ǹR�?rm$�� B�X��l?_ЯE��9�(�)�Z�ܣB����K�$����A,"�_A(��1w)b��U�>s�G�SS'pϡ�1�%� �w�$�O�j���1��p�*4�=���-zu��iBK��(��Tm�U�;�����6�S>����sliȀƅ�s|:�}��q��Dܱܭ�V��7���f+�e��T�q.�0�6P��E<�c���tc�����f�����x6Y�5�E	5P����M9I��9�b��Z�wal(�lipb>�q��t+M7��D}&���ǀ(}��l���v��춐���:�G�YԈ7n�� ���VJk�V�q�/F�d2��}�V5"*> ������.� ��
o�Cd~���� �����%�ېn�" �|��0%5���Nc|�7�� ��0�?&"�H�-�7II}t�R,	�y�gY�3<g�������O���+�e����!Wx�a c&��J���r���
���NݮÒ�@�,�N{�h������AU�j�aX����Cm��_9$���_P�Ey�H܃(f�g��l'@S=A4la�4���9�f��)o���R�q��X"��>��S��@[ui��
�./Pn�F�]�䇄O���
�"�(��\�F����i�W+�}N����E=������zf�W k�^�o-:�C��M��B��xE�!��ǘ���r*I#"��{`"�G�����E3���?��B�oA;���T�Bo�����~A�����$^���k�zC��|��u�J1�$�[z�0|qq��-����ϗ�yT�����E��r�t�C���x_�UJn�����c7��Q73���j��`C�|,����T���d��%�g�'#�����_e�qd�	�/:8���%�:�%����iW����䲪��#?\��D�ҕTaY-�p=��^ed�șiۗ��Pe��X8g�UMЈ������5�+ >��'��9v[�	��~'B���ʣ��F�CAi�&�V�2[���R�L��^������o����J����� ml��T��j9|gr9q&�6� ����pbJ�j@؅�\F|�
�B��,E2��ǿ����:�S�"0�'C���3�e���x1�� g*���%Yl�j��z�0"2[C��{QXv�~y�$�<ȉì�����)�
f"��f��p�~��W��=�х}�^�`���t�В4���/롧��ƞ2S��cm0c���=�->
���4���䃗8
}u�e\OK��T���6E&Xթ�R�^}2��[+���hJb�����~�%��+,�K�ۼZ�GV�e�"�o�]�^ʣh�'7��n|����Z����J�m]?����|���Ŝʦ K,���:�`{B�sq����k ��%�\�R��:g.�$����j��:1�-⻜.`��0��9~��\[H��r�!�i�v�RW5n�Dj!���(�l&3�� �
zR�TF��}�B�u�g(�赴�^��7��u��*1�>=J �u#
���<��kE�Z�t�\rO;\8���(8�Vբ2����^l�k>m���Z�};؇�j5j�ߴ�R�˒B��s��-g��'�}��g��x��WCLXAe��G�SkР�&�z��	����WB$F�!o7�V3E�gU8B�z�;�/
U��������[[��TW���~T�����s>4�IƋ�H��TmK��aʠ
�K�j�u����jf��9�O���n<��Vԛ���N�h�lg@�C�q:�[���ei2.mU�~*�����D�\��V�w�w���iͧ��k��1�+-�j�J�MSI6;-÷�x���vYd��'/�@�Y���
�r�cI�� �Sk*��,-���TO�	B�R�,m���&����{PQ30�̤N�7��a��O�R��1W�]���g`����m���Ji�=�8Y
x[E�.����H�^���HH�OW�e�����y��<�.��Dn���.PU���fG�*7~�U��Q��o�{{��F7�+�aA��T�±y-������C����� vU���IG�)��-iQF����4��.b2r<{pԿ�՛:2��߹"@1��h��}�]�z4h��_0���5i��̳��>V��j��q65�-iV��s�&N&�SyZ�ַ�@�C[��QE�T��D��������.w�4��R<�Qqo���6��:���he4�y>HFu�XK�#��Z���?/�$u��4��������oX�P<���. kM*[����V���A�^�CJ�,��#��f�e8�7.�q��'9�@��P��k
�ş��'o���I,��`��#��O��djW�w�d[EeQ�B�X l��
�w��ZQ0�*9Ћ��5W˗l�G#�c��:A����I�ٹ��/�!: jјQM#��#޵r'8������6w�X�zz(ʀtv4��p����5�]�Tjb����mxy����R[�h]���'z�A(��pC�4�pPzL�0�.dW?��@'G���]&�����D$jws8��QF!K����S:w��
g�\:� ֤�A��M=�k�M���<���Qa$����k�}���3$�&ɼܠL.p7iCsu�F60��1s�!Be��6-x-���nӾ�\ �������)���!L�[�+���-!����ݧ�4�5p��x|���K��C"����V�y��z��O0x� ��\�'�2��b�ֵ��$O�?�	/a�n��<v��Y���FS�X��ts����h�����,(7B��'�J��A�VH(q1��#>j[=�?q12)B�1�#��c�?D�ip5��ONt�2c�)�lU1oT~ p3׾Cb���ب�p��o� ��Q�l/ˣN�u��(����MT6�&d����eQ�	~�0>O�9o@�[Nw��\�v����f� ����˺��U6[�0F4��|$`�z�c�%U	�3���p��.�}�Ӟ��:bV_�8�n-�M�[w�<g�I�cC�o�b��'�ϧ,fJ�����mS${^v��ٻ�򨏵۷R���7�����c.�mӇb
7�A ����F���,	�d:�^��] �<D'3QO�|�|(*�Aut5��9tBF�J/�r�ڝ�?	����хw�>�}�� H��~� q���ڰ��>T�����y����=���7s����T�l����(�zod���u����~�ۛ��q{)^�)CL���.��><|d���D���Q�}�����r�74��i�2�P��	�(���,� �`��da��d���	����EQ�cB�ERd|�"_x�<�r*Ֆ|����C�.��<���f�6��s��(�n���!S���W�Z�;�E ������:�����O�!��05q����Y@��Cղ�=�|���d�sQ,�O'a�C&��L�=�D�~V!c����1��Nd��`lp
`�-���|��
���`VP)���$����I��C�K�%�h��;xS��/��{�f�@u8!��(���1kZ#y��m��l�Pi�$kM�	.d�=Ԑ�|���y�
���&ME2�	�}w[�����y�s���d�3]���Ѯ��¥}F�t�������`��D��Wɂ�����R��qX���f�mB���%M��1^��=�;r"D[���|�މ���W^撁Z&�߉�hdK�%�ve����@NMw�q�C���=�$gv����,�X��R@��9�����@�����	��b�Ṵ(�Y̌ȴ�}M�^����,�<�yT,/��������`_힎��Ș]
L+��ޙ[#��vl��c� @��?fyS�Bl�yP��(O��װ�/��w�=��3u
]����D����2�)�sw�|��i?b�(m��ke��[r�){n�+YI4<�y�H{�%�I~^�������3�Pj�b��Ŝ(`6Xxt+4���RԼ98j��[JւQ���@�q��-�R �)k�1s��2-]��$�&iI��X����e.s,ΒP@`lDHz/��>���e��u3?�%�:�jz�X�zR�C������_���D�а9`�����ѕ6�-�_po�h�<���5�R�Wt.���/ƛ�z~1ӎTCX�	Щ�f���5��M �')E�����G��r�gn���><Z�X��]D������u&gw*gk ���ge�I5b�O�M�Ϝ^�C8%k�� "=����U�jb��?s��"��	$���;���?%(��~[�֗RK��u:/b��V[,�j��z1m�E�����A�c�)WU�|��d�=f�Z��SkSꈒ�-7��%� '|����=�x��9ϭ��\|m@���*X�5���Zl�n50�\W�"KL]_m��;��A'�ꛆS�ã���BI~���{#cL����U�r�&�2�J��^��#A�O]kP��1'$+S��4���w��Ċ��	� �a�~���K����2s`�����)	��7�I7S9���lx�4����;M!Q����+m�P����GHz��/f#�]��Pd��;`G�&R�QΡ��[�+����嫻b�A_�.�_V,6ֳ6��`U�9<�����a��Jgx�L5t��}'C���c��6�C�"=K�ڍ+ϭ��`��2`���?n�SkA���F��Q�M�BM6*��/�D偂�+�OI�D!"T�؜�¯�e@T!�D�P*�}�ͧ��bvV�R?z�W��}�B^ʈQ��έd��x�<�p��0�-�=)�vl9������܊�s�RH�o9@�`ފ_�����|�F!go���D�]VE��%���͎�P,Y�����]��Q+���v7D�)���A���I�
�. �^�|�ﰆ*�mO���z����عM ���y@���6i�RŔx5Sc�����B�b?ynf&t.���8��Í�#��I]���ʢ���x��!�[�����@b�zjU��a���:��v�\�bt�2�<���_�o���gՒ�_t��h�\�tո����/Ǐ�;��t�"�YVu�)��� An�;�?�>��F�̦��k�q`|�Ec�N�A�X�˰;�jK�1��֭R"�^=-��i:z����1�9�ga���G�g�qX@��m�ѭ��H�N���c�8����4���1�M�%	C���O�����ܝ�F�󙯞M�G/��_/�w��h� �['�e�6�$;XKz�˼cp�e3�G�#�܁��%S�� EKr��n���}�L�I�ODʶ�*�S*l:�hcy�~�^)υ>��/�
A^ohS-�� ��1�����������կ	���m��õ�{�1�L0L�Դ�	�]�����t�_k۾�7Y;jN�=�zh�e�T-���9S�Y�?�l���Ђ��jH�볔~��`�9 ��׵���ᓶV}HJ�hq�g�$>,��Lm���E_�,2T��րw9	=���l��~��'`o�6��iՎPв��6/�3ꞧ�=<�_�S��15k
��&[��P <�4�S��x�s� :Wц��td����'�Ć�Q.��Q����/�Y�^;Ks`i�G������|��i��x^P�r^m�*P!)~�Ku�����"�j��F=�pʥ��a��a{�"Ø�F Q9�����;vrVr�V������R,��M���&� s���e]-��Gi!����e�ou�T�31���8lQ�HAnI(�L�#����� �}�y�w��6�K�^4^f�!c�l�n�Э�ח�H��0��-V��'jgP!�M*m]�,Y��&���x`&�]R{�7��?2�;�J q�&P��	�f�]M��h���Qz���XSJ����k��G{�]c�~2��,���.D�"�1�����Ȁ��cz; ��+w�ߓM|��I�Ry��{����x��?���R�]m?Wؼ�yE�s��5ߒ�԰aV0����+�ƥ��f˂D��-�;�����>�rQ����US0�V�DJ�9Q�/Fш���l	 l`os��u�Y���+~�I���⸎Q�2�~��t�;��@=�Ox~�����Hpg6n6jV��Gu��1RY�MC����&���.��偫J���n{S��*�9����g�md��PW�K�����Y��|����9��"v�p���K�P��]�;����L��(�Ӆ����J�Ѿ�/W�o�B�Ѹ��Aܺ(�,iN�{�}���̓��aaO)��\����vk-y}
��m>�f��n�@w�����⡯QS\�W�T�}�O��wG�T�:Ol�B���T�@*WU͕��U��(��&�"|I~��+X�V�_�Z8�C�~	9sM��󱟚�k�GZ�uy����z�t�*�`�2 �!�Xx݈����<~j��^�g*�%`�
]=��K���:d��K|D�P�z��p����(.�騱U0
�D^8�-�xۻ����I�(G�@ qE��r�s��ś��t�N�Y��C�d2b����z
�W��c Z�ڍ�o�oP8�
�Q^3U݇	b����?,WTN'�2���¾�P����H�2�2��u��6����(��b�8��J�H�3׺\Z�R��ESpdFB����u�b��E'�����q�����w�su�o��>c����U6ZF����Jd$7/T�e�l�X�k̢��ab��8��r�*���}H�&���u�� �S t���2P.�v���'+��89�"��Rg�s�
Q F5�$v��@ϝ�B�ck�v5���$��|ۜ&?1ʑ��ҕ6��^�{��2X�3��v���{��&9;p���[�W%���"��xa&b����͞�c�%6�F����6���T����%�$v��O��>�)0��k�n->P�qE���|�lĨ������K���4���p��	��=&��)�uQ0oJ�Hl�X?��$���f%��� �FU���6���KuU��`�q����o�Vո�7�	^cM���:z��1w�&�*
��$��82�P�F��ޜ/8��	�`�b��7�ۖ����o�b�ү��Jx9��QK�yP8��G+�yM�"�:�V��D��.K�����L�cD;�X�L�e����[��r;��=�Hk�k"����������2�� �`gfi?R�s;k��S�
�sa'v�sJ�,����s(��Ɉ8*7.iq��ed�78�[���J܁�&p�0M,��+�8��Y6uU�}�����I������F~�Ɉ��0�m�'c_�Ӎϩ��;U\p�J~-��׳�ַ��`{*z� s��O5�e�^��`=Q��K���;&v��w_�x��L`ϬҤ*�����;��W�n/�lK�fbI�i��d��sޥ�R	8]�)WJ�)"� x��ݒ��e2�3j`Mb�J �*]GjxC�A�?c��ۯf+-
HJ;8�@`�7Z��ߍ�
[��ZT�1Yߠ�qo8׼���\��� ����fB��w�&N&>R�;u��vW��$#�h��`��a���l�r���N ���<���㶂O��
��3�&�ȅ.�Rp^a!��$��q�N�zGT�����Kr?�߬�s:&CL��Ҿ,	j����[�$��
�el7�����䱸�	��fW��p;��}�ڈ�d�	U��Q���^~hD-͑�Z)��0���l[b�S�!Y�P�������u[��2��7i�����k�H\�,o��}1�u��m(Xqh���纀�������z`��Z<���3�\�	���I�����R�%)=�Tk0٬�"#a����IA<���y�\���X�����(�gp�WT�eZ0G�U ��+���s��&�A���̣,<��x��F���
R��fd\-*�3*���a�˻��#|�q<���IyRaxt��!˷m+���a`��0�T�����SR��2�U��5��a3�
5��F���D.��}Ԩ�݇9���z8KIz��T��]$����2|�#�����OԼm�/�d�Q�*�������,������h>����>C&::k=�m^Y=mY�*�����m�=�zޯCx�=|��I1�p���N��8� �t��ƻ��ו��^���/�����ҵ���DF���/ӈ�iF�x��8��7���ߟs�����A{&U�h����L���^9�D��]��Q��y��H��r�*���[��ewbyf^<~"�Ś��Z*<�%�!Gh&�ސ�?��cL����o��M�꿵/Mp��:�bxZtE��>�}[��
��>[܇W#EO]L�a�4゠y�"�L^΍�_��s-&m.�6�k�wY��4���T�5m[��c@w��)��9<�TmD��&���2��z���҆a����<Z���uϾ�G.yJ�O�B����4�kC�J��Y�n��7���g=�Nn|}�o��Z;s�s��"��&�%���0��p5g�;�z��)�_���I��3�Z��k�z)�2�}�{n�	o_ ag2ZI�wV!�>��*��1/A$qb�I�<����!9��a3v��m>ZW��4���
a�H��̮�$b�"2��+:GA6�نm����;Z���!�7@8춇^��c�)��vݵ�ۦ�Q��k�ϥ0{эU��h�H�쁿�  h���$M �%��=ti<7��*�B�U�E狥/��	��?۾��Ȫ��v��J�
��l�9��2@�������}�:������F��v/2���%��/�~��F!���q�&�HvW��� �dZ��?�����-�o+�����8a3<(��ҽ��/�6�r�U��4��ï��o�z�cQX�Gw�����=9T��8t�Y�H�֭����G{)�ӔA�l*O���x�~����H���I��e4��>D�XpTG��S���'uB�t��2�s���<a��8�֧^� ��+��Jm���Q#�	�ae�&�1q�ż�*�0�n�˸ӈ�[���*˴�Htzf�@t�#�"�]P���#��s�D%5[�&����D;�BY�r5Zq[8�s�	��Wc�O<�[J�-EV%G[n�U��m�Ɓ3��Qw�$�R(��#}.�,7s$�G�Ud{)k�8X�8�P��ʻ2(���x˗���;րv ��v�g[:�l�;��0d�VTN�t��U�9�tXu�.e`��)?���ϑ3P=9v����̄��V�Qwz4�ү�lY�^�������X����p�M��X���?*]gi�0���Ӳ?m�+pa�q��0�g�kY�Z�����5!����SU��aW	0�������V����8j���-闂>oD�J�3\8VB��,���wDM�Z�1.�B�H�X }D�É�y������D�6"�LN�9 h��z���m�'�z�vW!��w�Y������:=��v$}���d=S��i���<on9eGHn��=�l��r%��� <��1�샰��Ü�)Tq�)���C�}w`��g������E^��y+�;G)��4�cC&k�� _bE�R��7>��α�5
Y��`��L��c+Ur�a+)1�7h3�����Gy�\J�G��o���� �<��#���N��I���j�!�Y�|��gku�_�(7w�ڡ�6����l����nM�w�����4Ҳ�UW"�/�6�!��B9��KKt,-d����[�N˕�b���U��.�/YO��`�*}���|�teZ]U�jʢW%�x�Nm�&��-:P�:�����3klp#�w��V��^��B�־Xe3�E}�H�#L�C8�Z'g�+{��5�7ؑ�o@:�a`D�����;��v������;�$���v��`熎�do���bd��Ow����o���b�sUQ��S�Y���4%��Vx���&#�����EO��49\�{ �'4��rl!Ow\�0tO���2�l�+8o�Wz��Kc�p'�|��E������5�x��a�q\���v��=�i4�>e�+�^��ޡ�<ę U �Xn@Dt�x�6�?�0�ֆo��(�6(�M*������_�c��HlD�%�n��LkX2�	.ږ�^s����8��pᏺ��?~glxVsnn5������5�OVo��dXs�C��<��F��YT.�<�^�hƏŋ	�`ܣ���rXf�{G�&��7h��m��4����������C���g=�<(Q_,�&ᨇM���ѣ$��1�A��`Z9�����.�����b^�9~7U:���������V�Uɩ�lK|�.�[s��@^�s���\t+1<@�J_�x�� ��w	/�^��Hv���'c�fS�c���q��s~�����>�F��~Ō\{tJ/P��K��o2a�f�RǷ�<�@���L%^-D}��B�9����1�y��":�m3pnN�CT.vd�����k��@����g�M�X��J�8�����(�h}&'+gD��H��@�-dʷ�# %���JyfZƃ"דT���ٳ����ZV����;��p�=�iӌ�������ý��e�W�2M߆Xte聆~�䵷q�r����`�,��{��-W�W��#�o4��׭3�x������`W����� z� ;a����M@HӉ"��8���H���`c��k�e��(�G�mU�f�p�����˦�ağ`�y�p�F8��&�Ʀf��0LҀ���x9���`���ly�_�l�A~�a۳(tk�!��<#���|����9�g���]��_c�AQ1�g`��s]�2��|ԩ���EAE&Ʉi�	N��a�Ӏt���`]R% ����zz�-��J*ȟ����
d���W�`�`ѐO��s��	�t"���2��nK]V�Hc;���_2�y8�>����h�@��@j�/r�u����kt�n,���ƨ��P��bvm�1�,HoDǪ�>�u�*�F���{Ӕ�x,��K�p���"�Xr�#bL��B��:��DH�Ŀ�o�4w:I����T�l�9