module nodes (restart, clk, audio_out, sw);
	output wire signed [15:0] audio_out;
	input clk, restart;
	input [17:0] sw;


	wire signed[17:0] vwire_0_0;
	reg signed[17:0] vreg_0_0;
	node n0_0(.left(vreg_1_0), .right(vreg_1_0), .up(vreg_0_1), .down(vreg_0_1), .clk(clk), .reset(restart), .resetval(18'b001010001011111010), .value(vwire_0_0), .sw(sw));
	wire signed[17:0] vwire_0_1;
	reg signed[17:0] vreg_0_1;
	node n0_1(.left(vreg_1_1), .right(vreg_1_1), .up(vreg_0_2), .down(vreg_0_0), .clk(clk), .reset(restart), .resetval(18'b000110001011011001), .value(vwire_0_1), .sw(sw));
	wire signed[17:0] vwire_0_2;
	reg signed[17:0] vreg_0_2;
	node n0_2(.left(vreg_1_2), .right(vreg_1_2), .up(vreg_0_3), .down(vreg_0_1), .clk(clk), .reset(restart), .resetval(18'b000001011000001110), .value(vwire_0_2), .sw(sw));
	wire signed[17:0] vwire_0_3;
	reg signed[17:0] vreg_0_3;
	node n0_3(.left(vreg_1_3), .right(vreg_1_3), .up(vreg_0_4), .down(vreg_0_2), .clk(clk), .reset(restart), .resetval(18'b000000000111001111), .value(vwire_0_3), .sw(sw));
	wire signed[17:0] vwire_0_4;
	reg signed[17:0] vreg_0_4;
	node n0_4(.left(vreg_1_4), .right(vreg_1_4), .up(vreg_0_5), .down(vreg_0_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_4), .sw(sw));
	wire signed[17:0] vwire_0_5;
	reg signed[17:0] vreg_0_5;
	node n0_5(.left(vreg_1_5), .right(vreg_1_5), .up(vreg_0_6), .down(vreg_0_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_5), .sw(sw));
	wire signed[17:0] vwire_0_6;
	reg signed[17:0] vreg_0_6;
	node n0_6(.left(vreg_1_6), .right(vreg_1_6), .up(vreg_0_7), .down(vreg_0_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_6), .sw(sw));
	wire signed[17:0] vwire_0_7;
	reg signed[17:0] vreg_0_7;
	node n0_7(.left(vreg_1_7), .right(vreg_1_7), .up(vreg_0_8), .down(vreg_0_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_7), .sw(sw));
	wire signed[17:0] vwire_0_8;
	reg signed[17:0] vreg_0_8;
	node n0_8(.left(vreg_1_8), .right(vreg_1_8), .up(vreg_0_9), .down(vreg_0_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_8), .sw(sw));
	wire signed[17:0] vwire_0_9;
	reg signed[17:0] vreg_0_9;
	node n0_9(.left(vreg_1_9), .right(vreg_1_9), .up(vreg_0_10), .down(vreg_0_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_9), .sw(sw));
	wire signed[17:0] vwire_0_10;
	reg signed[17:0] vreg_0_10;
	node n0_10(.left(vreg_1_10), .right(vreg_1_10), .up(vreg_0_11), .down(vreg_0_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_10), .sw(sw));
	wire signed[17:0] vwire_0_11;
	reg signed[17:0] vreg_0_11;
	node n0_11(.left(vreg_1_11), .right(vreg_1_11), .up(vreg_0_12), .down(vreg_0_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_11), .sw(sw));
	wire signed[17:0] vwire_0_12;
	reg signed[17:0] vreg_0_12;
	node n0_12(.left(vreg_1_12), .right(vreg_1_12), .up(vreg_0_13), .down(vreg_0_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_12), .sw(sw));
	wire signed[17:0] vwire_0_13;
	reg signed[17:0] vreg_0_13;
	node n0_13(.left(vreg_1_13), .right(vreg_1_13), .up(vreg_0_14), .down(vreg_0_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_13), .sw(sw));
	wire signed[17:0] vwire_0_14;
	reg signed[17:0] vreg_0_14;
	node n0_14(.left(vreg_1_14), .right(vreg_1_14), .up(vreg_0_15), .down(vreg_0_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_14), .sw(sw));
	wire signed[17:0] vwire_0_15;
	reg signed[17:0] vreg_0_15;
	node n0_15(.left(vreg_1_15), .right(vreg_1_15), .up(vreg_0_16), .down(vreg_0_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_15), .sw(sw));
	wire signed[17:0] vwire_0_16;
	reg signed[17:0] vreg_0_16;
	node n0_16(.left(vreg_1_16), .right(vreg_1_16), .up(vreg_0_17), .down(vreg_0_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_16), .sw(sw));
	wire signed[17:0] vwire_0_17;
	reg signed[17:0] vreg_0_17;
	node n0_17(.left(vreg_1_17), .right(vreg_1_17), .up(vreg_0_18), .down(vreg_0_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_17), .sw(sw));
	wire signed[17:0] vwire_0_18;
	reg signed[17:0] vreg_0_18;
	node n0_18(.left(vreg_1_18), .right(vreg_1_18), .up(vreg_0_19), .down(vreg_0_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_18), .sw(sw));
	wire signed[17:0] vwire_0_19;
	reg signed[17:0] vreg_0_19;
	node n0_19(.left(vreg_1_19), .right(vreg_1_19), .up(vreg_0_20), .down(vreg_0_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_19), .sw(sw));
	wire signed[17:0] vwire_0_20;
	reg signed[17:0] vreg_0_20;
	node n0_20(.left(vreg_1_20), .right(vreg_1_20), .up(vreg_0_21), .down(vreg_0_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_20), .sw(sw));
	wire signed[17:0] vwire_0_21;
	reg signed[17:0] vreg_0_21;
	node n0_21(.left(vreg_1_21), .right(vreg_1_21), .up(vreg_0_22), .down(vreg_0_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_21), .sw(sw));
	wire signed[17:0] vwire_0_22;
	reg signed[17:0] vreg_0_22;
	node n0_22(.left(vreg_1_22), .right(vreg_1_22), .up(vreg_0_23), .down(vreg_0_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_22), .sw(sw));
	wire signed[17:0] vwire_0_23;
	reg signed[17:0] vreg_0_23;
	node n0_23(.left(vreg_1_23), .right(vreg_1_23), .up(vreg_0_24), .down(vreg_0_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_23), .sw(sw));
	wire signed[17:0] vwire_0_24;
	reg signed[17:0] vreg_0_24;
	node n0_24(.left(vreg_1_24), .right(vreg_1_24), .up(vreg_0_25), .down(vreg_0_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_24), .sw(sw));
	wire signed[17:0] vwire_0_25;
	reg signed[17:0] vreg_0_25;
	node n0_25(.left(vreg_1_25), .right(vreg_1_25), .up(vreg_0_26), .down(vreg_0_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_25), .sw(sw));
	wire signed[17:0] vwire_0_26;
	reg signed[17:0] vreg_0_26;
	node n0_26(.left(vreg_1_26), .right(vreg_1_26), .up(vreg_0_27), .down(vreg_0_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_26), .sw(sw));
	wire signed[17:0] vwire_0_27;
	reg signed[17:0] vreg_0_27;
	node n0_27(.left(vreg_1_27), .right(vreg_1_27), .up(vreg_0_28), .down(vreg_0_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_27), .sw(sw));
	wire signed[17:0] vwire_0_28;
	reg signed[17:0] vreg_0_28;
	node n0_28(.left(vreg_1_28), .right(vreg_1_28), .up(vreg_0_29), .down(vreg_0_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_28), .sw(sw));
	wire signed[17:0] vwire_0_29;
	reg signed[17:0] vreg_0_29;
	node n0_29(.left(vreg_1_29), .right(vreg_1_29), .up(vreg_0_30), .down(vreg_0_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_29), .sw(sw));
	wire signed[17:0] vwire_0_30;
	reg signed[17:0] vreg_0_30;
	node n0_30(.left(vreg_1_30), .right(vreg_1_30), .up(vreg_0_31), .down(vreg_0_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_30), .sw(sw));
	wire signed[17:0] vwire_0_31;
	reg signed[17:0] vreg_0_31;
	node n0_31(.left(vreg_1_31), .right(vreg_1_31), .up(vreg_0_32), .down(vreg_0_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_31), .sw(sw));
	wire signed[17:0] vwire_0_32;
	reg signed[17:0] vreg_0_32;
	node n0_32(.left(vreg_1_32), .right(vreg_1_32), .up(vreg_0_33), .down(vreg_0_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_32), .sw(sw));
	wire signed[17:0] vwire_0_33;
	reg signed[17:0] vreg_0_33;
	node n0_33(.left(vreg_1_33), .right(vreg_1_33), .up(vreg_0_34), .down(vreg_0_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_33), .sw(sw));
	wire signed[17:0] vwire_0_34;
	reg signed[17:0] vreg_0_34;
	node n0_34(.left(vreg_1_34), .right(vreg_1_34), .up(vreg_0_35), .down(vreg_0_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_34), .sw(sw));
	wire signed[17:0] vwire_0_35;
	reg signed[17:0] vreg_0_35;
	node n0_35(.left(vreg_1_35), .right(vreg_1_35), .up(vreg_0_36), .down(vreg_0_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_35), .sw(sw));
	wire signed[17:0] vwire_0_36;
	reg signed[17:0] vreg_0_36;
	node n0_36(.left(vreg_1_36), .right(vreg_1_36), .up(vreg_0_37), .down(vreg_0_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_36), .sw(sw));
	wire signed[17:0] vwire_0_37;
	reg signed[17:0] vreg_0_37;
	node n0_37(.left(vreg_1_37), .right(vreg_1_37), .up(vreg_0_38), .down(vreg_0_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_37), .sw(sw));
	wire signed[17:0] vwire_0_38;
	reg signed[17:0] vreg_0_38;
	node n0_38(.left(vreg_1_38), .right(vreg_1_38), .up(vreg_0_39), .down(vreg_0_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_38), .sw(sw));
	wire signed[17:0] vwire_0_39;
	reg signed[17:0] vreg_0_39;
	node n0_39(.left(vreg_1_39), .right(vreg_1_39), .up(vreg_0_40), .down(vreg_0_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_39), .sw(sw));
	wire signed[17:0] vwire_0_40;
	reg signed[17:0] vreg_0_40;
	node n0_40(.left(vreg_1_40), .right(vreg_1_40), .up(vreg_0_41), .down(vreg_0_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_40), .sw(sw));
	wire signed[17:0] vwire_0_41;
	reg signed[17:0] vreg_0_41;
	node n0_41(.left(vreg_1_41), .right(vreg_1_41), .up(vreg_0_42), .down(vreg_0_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_41), .sw(sw));
	wire signed[17:0] vwire_0_42;
	reg signed[17:0] vreg_0_42;
	node n0_42(.left(vreg_1_42), .right(vreg_1_42), .up(vreg_0_43), .down(vreg_0_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_42), .sw(sw));
	wire signed[17:0] vwire_0_43;
	reg signed[17:0] vreg_0_43;
	node n0_43(.left(vreg_1_43), .right(vreg_1_43), .up(vreg_0_44), .down(vreg_0_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_43), .sw(sw));
	wire signed[17:0] vwire_0_44;
	reg signed[17:0] vreg_0_44;
	node n0_44(.left(vreg_1_44), .right(vreg_1_44), .up(vreg_0_45), .down(vreg_0_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_44), .sw(sw));
	wire signed[17:0] vwire_0_45;
	reg signed[17:0] vreg_0_45;
	node n0_45(.left(vreg_1_45), .right(vreg_1_45), .up(vreg_0_46), .down(vreg_0_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_45), .sw(sw));
	wire signed[17:0] vwire_0_46;
	reg signed[17:0] vreg_0_46;
	node n0_46(.left(vreg_1_46), .right(vreg_1_46), .up(vreg_0_47), .down(vreg_0_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_46), .sw(sw));
	wire signed[17:0] vwire_0_47;
	reg signed[17:0] vreg_0_47;
	node n0_47(.left(vreg_1_47), .right(vreg_1_47), .up(vreg_0_48), .down(vreg_0_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_47), .sw(sw));
	wire signed[17:0] vwire_0_48;
	reg signed[17:0] vreg_0_48;
	node n0_48(.left(vreg_1_48), .right(vreg_1_48), .up(vreg_0_49), .down(vreg_0_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_48), .sw(sw));
	wire signed[17:0] vwire_0_49;
	reg signed[17:0] vreg_0_49;
	node n0_49(.left(vreg_1_49), .right(vreg_1_49), .up(18'b0), .down(vreg_0_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_49), .sw(sw));
	wire signed[17:0] vwire_1_0;
	reg signed[17:0] vreg_1_0;
	node n1_0(.left(vreg_0_0), .right(vreg_2_0), .up(vreg_1_1), .down(vreg_1_1), .clk(clk), .reset(restart), .resetval(18'b000110001011011001), .value(vwire_1_0), .sw(sw));
	wire signed[17:0] vwire_1_1;
	reg signed[17:0] vreg_1_1;
	node n1_1(.left(vreg_0_1), .right(vreg_2_1), .up(vreg_1_2), .down(vreg_1_0), .clk(clk), .reset(restart), .resetval(18'b000011101111110100), .value(vwire_1_1), .sw(sw));
	wire signed[17:0] vwire_1_2;
	reg signed[17:0] vreg_1_2;
	node n1_2(.left(vreg_0_2), .right(vreg_2_2), .up(vreg_1_3), .down(vreg_1_1), .clk(clk), .reset(restart), .resetval(18'b000000110101100001), .value(vwire_1_2), .sw(sw));
	wire signed[17:0] vwire_1_3;
	reg signed[17:0] vreg_1_3;
	node n1_3(.left(vreg_0_3), .right(vreg_2_3), .up(vreg_1_4), .down(vreg_1_2), .clk(clk), .reset(restart), .resetval(18'b000000000100011001), .value(vwire_1_3), .sw(sw));
	wire signed[17:0] vwire_1_4;
	reg signed[17:0] vreg_1_4;
	node n1_4(.left(vreg_0_4), .right(vreg_2_4), .up(vreg_1_5), .down(vreg_1_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_4), .sw(sw));
	wire signed[17:0] vwire_1_5;
	reg signed[17:0] vreg_1_5;
	node n1_5(.left(vreg_0_5), .right(vreg_2_5), .up(vreg_1_6), .down(vreg_1_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_5), .sw(sw));
	wire signed[17:0] vwire_1_6;
	reg signed[17:0] vreg_1_6;
	node n1_6(.left(vreg_0_6), .right(vreg_2_6), .up(vreg_1_7), .down(vreg_1_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_6), .sw(sw));
	wire signed[17:0] vwire_1_7;
	reg signed[17:0] vreg_1_7;
	node n1_7(.left(vreg_0_7), .right(vreg_2_7), .up(vreg_1_8), .down(vreg_1_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_7), .sw(sw));
	wire signed[17:0] vwire_1_8;
	reg signed[17:0] vreg_1_8;
	node n1_8(.left(vreg_0_8), .right(vreg_2_8), .up(vreg_1_9), .down(vreg_1_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_8), .sw(sw));
	wire signed[17:0] vwire_1_9;
	reg signed[17:0] vreg_1_9;
	node n1_9(.left(vreg_0_9), .right(vreg_2_9), .up(vreg_1_10), .down(vreg_1_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_9), .sw(sw));
	wire signed[17:0] vwire_1_10;
	reg signed[17:0] vreg_1_10;
	node n1_10(.left(vreg_0_10), .right(vreg_2_10), .up(vreg_1_11), .down(vreg_1_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_10), .sw(sw));
	wire signed[17:0] vwire_1_11;
	reg signed[17:0] vreg_1_11;
	node n1_11(.left(vreg_0_11), .right(vreg_2_11), .up(vreg_1_12), .down(vreg_1_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_11), .sw(sw));
	wire signed[17:0] vwire_1_12;
	reg signed[17:0] vreg_1_12;
	node n1_12(.left(vreg_0_12), .right(vreg_2_12), .up(vreg_1_13), .down(vreg_1_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_12), .sw(sw));
	wire signed[17:0] vwire_1_13;
	reg signed[17:0] vreg_1_13;
	node n1_13(.left(vreg_0_13), .right(vreg_2_13), .up(vreg_1_14), .down(vreg_1_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_13), .sw(sw));
	wire signed[17:0] vwire_1_14;
	reg signed[17:0] vreg_1_14;
	node n1_14(.left(vreg_0_14), .right(vreg_2_14), .up(vreg_1_15), .down(vreg_1_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_14), .sw(sw));
	wire signed[17:0] vwire_1_15;
	reg signed[17:0] vreg_1_15;
	node n1_15(.left(vreg_0_15), .right(vreg_2_15), .up(vreg_1_16), .down(vreg_1_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_15), .sw(sw));
	wire signed[17:0] vwire_1_16;
	reg signed[17:0] vreg_1_16;
	node n1_16(.left(vreg_0_16), .right(vreg_2_16), .up(vreg_1_17), .down(vreg_1_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_16), .sw(sw));
	wire signed[17:0] vwire_1_17;
	reg signed[17:0] vreg_1_17;
	node n1_17(.left(vreg_0_17), .right(vreg_2_17), .up(vreg_1_18), .down(vreg_1_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_17), .sw(sw));
	wire signed[17:0] vwire_1_18;
	reg signed[17:0] vreg_1_18;
	node n1_18(.left(vreg_0_18), .right(vreg_2_18), .up(vreg_1_19), .down(vreg_1_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_18), .sw(sw));
	wire signed[17:0] vwire_1_19;
	reg signed[17:0] vreg_1_19;
	node n1_19(.left(vreg_0_19), .right(vreg_2_19), .up(vreg_1_20), .down(vreg_1_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_19), .sw(sw));
	wire signed[17:0] vwire_1_20;
	reg signed[17:0] vreg_1_20;
	node n1_20(.left(vreg_0_20), .right(vreg_2_20), .up(vreg_1_21), .down(vreg_1_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_20), .sw(sw));
	wire signed[17:0] vwire_1_21;
	reg signed[17:0] vreg_1_21;
	node n1_21(.left(vreg_0_21), .right(vreg_2_21), .up(vreg_1_22), .down(vreg_1_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_21), .sw(sw));
	wire signed[17:0] vwire_1_22;
	reg signed[17:0] vreg_1_22;
	node n1_22(.left(vreg_0_22), .right(vreg_2_22), .up(vreg_1_23), .down(vreg_1_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_22), .sw(sw));
	wire signed[17:0] vwire_1_23;
	reg signed[17:0] vreg_1_23;
	node n1_23(.left(vreg_0_23), .right(vreg_2_23), .up(vreg_1_24), .down(vreg_1_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_23), .sw(sw));
	wire signed[17:0] vwire_1_24;
	reg signed[17:0] vreg_1_24;
	node n1_24(.left(vreg_0_24), .right(vreg_2_24), .up(vreg_1_25), .down(vreg_1_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_24), .sw(sw));
	wire signed[17:0] vwire_1_25;
	reg signed[17:0] vreg_1_25;
	node n1_25(.left(vreg_0_25), .right(vreg_2_25), .up(vreg_1_26), .down(vreg_1_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_25), .sw(sw));
	wire signed[17:0] vwire_1_26;
	reg signed[17:0] vreg_1_26;
	node n1_26(.left(vreg_0_26), .right(vreg_2_26), .up(vreg_1_27), .down(vreg_1_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_26), .sw(sw));
	wire signed[17:0] vwire_1_27;
	reg signed[17:0] vreg_1_27;
	node n1_27(.left(vreg_0_27), .right(vreg_2_27), .up(vreg_1_28), .down(vreg_1_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_27), .sw(sw));
	wire signed[17:0] vwire_1_28;
	reg signed[17:0] vreg_1_28;
	node n1_28(.left(vreg_0_28), .right(vreg_2_28), .up(vreg_1_29), .down(vreg_1_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_28), .sw(sw));
	wire signed[17:0] vwire_1_29;
	reg signed[17:0] vreg_1_29;
	node n1_29(.left(vreg_0_29), .right(vreg_2_29), .up(vreg_1_30), .down(vreg_1_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_29), .sw(sw));
	wire signed[17:0] vwire_1_30;
	reg signed[17:0] vreg_1_30;
	node n1_30(.left(vreg_0_30), .right(vreg_2_30), .up(vreg_1_31), .down(vreg_1_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_30), .sw(sw));
	wire signed[17:0] vwire_1_31;
	reg signed[17:0] vreg_1_31;
	node n1_31(.left(vreg_0_31), .right(vreg_2_31), .up(vreg_1_32), .down(vreg_1_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_31), .sw(sw));
	wire signed[17:0] vwire_1_32;
	reg signed[17:0] vreg_1_32;
	node n1_32(.left(vreg_0_32), .right(vreg_2_32), .up(vreg_1_33), .down(vreg_1_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_32), .sw(sw));
	wire signed[17:0] vwire_1_33;
	reg signed[17:0] vreg_1_33;
	node n1_33(.left(vreg_0_33), .right(vreg_2_33), .up(vreg_1_34), .down(vreg_1_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_33), .sw(sw));
	wire signed[17:0] vwire_1_34;
	reg signed[17:0] vreg_1_34;
	node n1_34(.left(vreg_0_34), .right(vreg_2_34), .up(vreg_1_35), .down(vreg_1_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_34), .sw(sw));
	wire signed[17:0] vwire_1_35;
	reg signed[17:0] vreg_1_35;
	node n1_35(.left(vreg_0_35), .right(vreg_2_35), .up(vreg_1_36), .down(vreg_1_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_35), .sw(sw));
	wire signed[17:0] vwire_1_36;
	reg signed[17:0] vreg_1_36;
	node n1_36(.left(vreg_0_36), .right(vreg_2_36), .up(vreg_1_37), .down(vreg_1_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_36), .sw(sw));
	wire signed[17:0] vwire_1_37;
	reg signed[17:0] vreg_1_37;
	node n1_37(.left(vreg_0_37), .right(vreg_2_37), .up(vreg_1_38), .down(vreg_1_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_37), .sw(sw));
	wire signed[17:0] vwire_1_38;
	reg signed[17:0] vreg_1_38;
	node n1_38(.left(vreg_0_38), .right(vreg_2_38), .up(vreg_1_39), .down(vreg_1_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_38), .sw(sw));
	wire signed[17:0] vwire_1_39;
	reg signed[17:0] vreg_1_39;
	node n1_39(.left(vreg_0_39), .right(vreg_2_39), .up(vreg_1_40), .down(vreg_1_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_39), .sw(sw));
	wire signed[17:0] vwire_1_40;
	reg signed[17:0] vreg_1_40;
	node n1_40(.left(vreg_0_40), .right(vreg_2_40), .up(vreg_1_41), .down(vreg_1_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_40), .sw(sw));
	wire signed[17:0] vwire_1_41;
	reg signed[17:0] vreg_1_41;
	node n1_41(.left(vreg_0_41), .right(vreg_2_41), .up(vreg_1_42), .down(vreg_1_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_41), .sw(sw));
	wire signed[17:0] vwire_1_42;
	reg signed[17:0] vreg_1_42;
	node n1_42(.left(vreg_0_42), .right(vreg_2_42), .up(vreg_1_43), .down(vreg_1_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_42), .sw(sw));
	wire signed[17:0] vwire_1_43;
	reg signed[17:0] vreg_1_43;
	node n1_43(.left(vreg_0_43), .right(vreg_2_43), .up(vreg_1_44), .down(vreg_1_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_43), .sw(sw));
	wire signed[17:0] vwire_1_44;
	reg signed[17:0] vreg_1_44;
	node n1_44(.left(vreg_0_44), .right(vreg_2_44), .up(vreg_1_45), .down(vreg_1_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_44), .sw(sw));
	wire signed[17:0] vwire_1_45;
	reg signed[17:0] vreg_1_45;
	node n1_45(.left(vreg_0_45), .right(vreg_2_45), .up(vreg_1_46), .down(vreg_1_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_45), .sw(sw));
	wire signed[17:0] vwire_1_46;
	reg signed[17:0] vreg_1_46;
	node n1_46(.left(vreg_0_46), .right(vreg_2_46), .up(vreg_1_47), .down(vreg_1_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_46), .sw(sw));
	wire signed[17:0] vwire_1_47;
	reg signed[17:0] vreg_1_47;
	node n1_47(.left(vreg_0_47), .right(vreg_2_47), .up(vreg_1_48), .down(vreg_1_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_47), .sw(sw));
	wire signed[17:0] vwire_1_48;
	reg signed[17:0] vreg_1_48;
	node n1_48(.left(vreg_0_48), .right(vreg_2_48), .up(vreg_1_49), .down(vreg_1_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_48), .sw(sw));
	wire signed[17:0] vwire_1_49;
	reg signed[17:0] vreg_1_49;
	node n1_49(.left(vreg_0_49), .right(vreg_2_49), .up(18'b0), .down(vreg_1_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_49), .sw(sw));
	wire signed[17:0] vwire_2_0;
	reg signed[17:0] vreg_2_0;
	node n2_0(.left(vreg_1_0), .right(vreg_3_0), .up(vreg_2_1), .down(vreg_2_1), .clk(clk), .reset(restart), .resetval(18'b000001011000001110), .value(vwire_2_0), .sw(sw));
	wire signed[17:0] vwire_2_1;
	reg signed[17:0] vreg_2_1;
	node n2_1(.left(vreg_1_1), .right(vreg_3_1), .up(vreg_2_2), .down(vreg_2_0), .clk(clk), .reset(restart), .resetval(18'b000000110101100001), .value(vwire_2_1), .sw(sw));
	wire signed[17:0] vwire_2_2;
	reg signed[17:0] vreg_2_2;
	node n2_2(.left(vreg_1_2), .right(vreg_3_2), .up(vreg_2_3), .down(vreg_2_1), .clk(clk), .reset(restart), .resetval(18'b000000001011111100), .value(vwire_2_2), .sw(sw));
	wire signed[17:0] vwire_2_3;
	reg signed[17:0] vreg_2_3;
	node n2_3(.left(vreg_1_3), .right(vreg_3_3), .up(vreg_2_4), .down(vreg_2_2), .clk(clk), .reset(restart), .resetval(18'b000000000000111111), .value(vwire_2_3), .sw(sw));
	wire signed[17:0] vwire_2_4;
	reg signed[17:0] vreg_2_4;
	node n2_4(.left(vreg_1_4), .right(vreg_3_4), .up(vreg_2_5), .down(vreg_2_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_4), .sw(sw));
	wire signed[17:0] vwire_2_5;
	reg signed[17:0] vreg_2_5;
	node n2_5(.left(vreg_1_5), .right(vreg_3_5), .up(vreg_2_6), .down(vreg_2_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_5), .sw(sw));
	wire signed[17:0] vwire_2_6;
	reg signed[17:0] vreg_2_6;
	node n2_6(.left(vreg_1_6), .right(vreg_3_6), .up(vreg_2_7), .down(vreg_2_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_6), .sw(sw));
	wire signed[17:0] vwire_2_7;
	reg signed[17:0] vreg_2_7;
	node n2_7(.left(vreg_1_7), .right(vreg_3_7), .up(vreg_2_8), .down(vreg_2_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_7), .sw(sw));
	wire signed[17:0] vwire_2_8;
	reg signed[17:0] vreg_2_8;
	node n2_8(.left(vreg_1_8), .right(vreg_3_8), .up(vreg_2_9), .down(vreg_2_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_8), .sw(sw));
	wire signed[17:0] vwire_2_9;
	reg signed[17:0] vreg_2_9;
	node n2_9(.left(vreg_1_9), .right(vreg_3_9), .up(vreg_2_10), .down(vreg_2_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_9), .sw(sw));
	wire signed[17:0] vwire_2_10;
	reg signed[17:0] vreg_2_10;
	node n2_10(.left(vreg_1_10), .right(vreg_3_10), .up(vreg_2_11), .down(vreg_2_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_10), .sw(sw));
	wire signed[17:0] vwire_2_11;
	reg signed[17:0] vreg_2_11;
	node n2_11(.left(vreg_1_11), .right(vreg_3_11), .up(vreg_2_12), .down(vreg_2_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_11), .sw(sw));
	wire signed[17:0] vwire_2_12;
	reg signed[17:0] vreg_2_12;
	node n2_12(.left(vreg_1_12), .right(vreg_3_12), .up(vreg_2_13), .down(vreg_2_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_12), .sw(sw));
	wire signed[17:0] vwire_2_13;
	reg signed[17:0] vreg_2_13;
	node n2_13(.left(vreg_1_13), .right(vreg_3_13), .up(vreg_2_14), .down(vreg_2_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_13), .sw(sw));
	wire signed[17:0] vwire_2_14;
	reg signed[17:0] vreg_2_14;
	node n2_14(.left(vreg_1_14), .right(vreg_3_14), .up(vreg_2_15), .down(vreg_2_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_14), .sw(sw));
	wire signed[17:0] vwire_2_15;
	reg signed[17:0] vreg_2_15;
	node n2_15(.left(vreg_1_15), .right(vreg_3_15), .up(vreg_2_16), .down(vreg_2_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_15), .sw(sw));
	wire signed[17:0] vwire_2_16;
	reg signed[17:0] vreg_2_16;
	node n2_16(.left(vreg_1_16), .right(vreg_3_16), .up(vreg_2_17), .down(vreg_2_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_16), .sw(sw));
	wire signed[17:0] vwire_2_17;
	reg signed[17:0] vreg_2_17;
	node n2_17(.left(vreg_1_17), .right(vreg_3_17), .up(vreg_2_18), .down(vreg_2_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_17), .sw(sw));
	wire signed[17:0] vwire_2_18;
	reg signed[17:0] vreg_2_18;
	node n2_18(.left(vreg_1_18), .right(vreg_3_18), .up(vreg_2_19), .down(vreg_2_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_18), .sw(sw));
	wire signed[17:0] vwire_2_19;
	reg signed[17:0] vreg_2_19;
	node n2_19(.left(vreg_1_19), .right(vreg_3_19), .up(vreg_2_20), .down(vreg_2_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_19), .sw(sw));
	wire signed[17:0] vwire_2_20;
	reg signed[17:0] vreg_2_20;
	node n2_20(.left(vreg_1_20), .right(vreg_3_20), .up(vreg_2_21), .down(vreg_2_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_20), .sw(sw));
	wire signed[17:0] vwire_2_21;
	reg signed[17:0] vreg_2_21;
	node n2_21(.left(vreg_1_21), .right(vreg_3_21), .up(vreg_2_22), .down(vreg_2_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_21), .sw(sw));
	wire signed[17:0] vwire_2_22;
	reg signed[17:0] vreg_2_22;
	node n2_22(.left(vreg_1_22), .right(vreg_3_22), .up(vreg_2_23), .down(vreg_2_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_22), .sw(sw));
	wire signed[17:0] vwire_2_23;
	reg signed[17:0] vreg_2_23;
	node n2_23(.left(vreg_1_23), .right(vreg_3_23), .up(vreg_2_24), .down(vreg_2_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_23), .sw(sw));
	wire signed[17:0] vwire_2_24;
	reg signed[17:0] vreg_2_24;
	node n2_24(.left(vreg_1_24), .right(vreg_3_24), .up(vreg_2_25), .down(vreg_2_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_24), .sw(sw));
	wire signed[17:0] vwire_2_25;
	reg signed[17:0] vreg_2_25;
	node n2_25(.left(vreg_1_25), .right(vreg_3_25), .up(vreg_2_26), .down(vreg_2_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_25), .sw(sw));
	wire signed[17:0] vwire_2_26;
	reg signed[17:0] vreg_2_26;
	node n2_26(.left(vreg_1_26), .right(vreg_3_26), .up(vreg_2_27), .down(vreg_2_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_26), .sw(sw));
	wire signed[17:0] vwire_2_27;
	reg signed[17:0] vreg_2_27;
	node n2_27(.left(vreg_1_27), .right(vreg_3_27), .up(vreg_2_28), .down(vreg_2_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_27), .sw(sw));
	wire signed[17:0] vwire_2_28;
	reg signed[17:0] vreg_2_28;
	node n2_28(.left(vreg_1_28), .right(vreg_3_28), .up(vreg_2_29), .down(vreg_2_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_28), .sw(sw));
	wire signed[17:0] vwire_2_29;
	reg signed[17:0] vreg_2_29;
	node n2_29(.left(vreg_1_29), .right(vreg_3_29), .up(vreg_2_30), .down(vreg_2_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_29), .sw(sw));
	wire signed[17:0] vwire_2_30;
	reg signed[17:0] vreg_2_30;
	node n2_30(.left(vreg_1_30), .right(vreg_3_30), .up(vreg_2_31), .down(vreg_2_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_30), .sw(sw));
	wire signed[17:0] vwire_2_31;
	reg signed[17:0] vreg_2_31;
	node n2_31(.left(vreg_1_31), .right(vreg_3_31), .up(vreg_2_32), .down(vreg_2_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_31), .sw(sw));
	wire signed[17:0] vwire_2_32;
	reg signed[17:0] vreg_2_32;
	node n2_32(.left(vreg_1_32), .right(vreg_3_32), .up(vreg_2_33), .down(vreg_2_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_32), .sw(sw));
	wire signed[17:0] vwire_2_33;
	reg signed[17:0] vreg_2_33;
	node n2_33(.left(vreg_1_33), .right(vreg_3_33), .up(vreg_2_34), .down(vreg_2_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_33), .sw(sw));
	wire signed[17:0] vwire_2_34;
	reg signed[17:0] vreg_2_34;
	node n2_34(.left(vreg_1_34), .right(vreg_3_34), .up(vreg_2_35), .down(vreg_2_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_34), .sw(sw));
	wire signed[17:0] vwire_2_35;
	reg signed[17:0] vreg_2_35;
	node n2_35(.left(vreg_1_35), .right(vreg_3_35), .up(vreg_2_36), .down(vreg_2_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_35), .sw(sw));
	wire signed[17:0] vwire_2_36;
	reg signed[17:0] vreg_2_36;
	node n2_36(.left(vreg_1_36), .right(vreg_3_36), .up(vreg_2_37), .down(vreg_2_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_36), .sw(sw));
	wire signed[17:0] vwire_2_37;
	reg signed[17:0] vreg_2_37;
	node n2_37(.left(vreg_1_37), .right(vreg_3_37), .up(vreg_2_38), .down(vreg_2_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_37), .sw(sw));
	wire signed[17:0] vwire_2_38;
	reg signed[17:0] vreg_2_38;
	node n2_38(.left(vreg_1_38), .right(vreg_3_38), .up(vreg_2_39), .down(vreg_2_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_38), .sw(sw));
	wire signed[17:0] vwire_2_39;
	reg signed[17:0] vreg_2_39;
	node n2_39(.left(vreg_1_39), .right(vreg_3_39), .up(vreg_2_40), .down(vreg_2_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_39), .sw(sw));
	wire signed[17:0] vwire_2_40;
	reg signed[17:0] vreg_2_40;
	node n2_40(.left(vreg_1_40), .right(vreg_3_40), .up(vreg_2_41), .down(vreg_2_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_40), .sw(sw));
	wire signed[17:0] vwire_2_41;
	reg signed[17:0] vreg_2_41;
	node n2_41(.left(vreg_1_41), .right(vreg_3_41), .up(vreg_2_42), .down(vreg_2_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_41), .sw(sw));
	wire signed[17:0] vwire_2_42;
	reg signed[17:0] vreg_2_42;
	node n2_42(.left(vreg_1_42), .right(vreg_3_42), .up(vreg_2_43), .down(vreg_2_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_42), .sw(sw));
	wire signed[17:0] vwire_2_43;
	reg signed[17:0] vreg_2_43;
	node n2_43(.left(vreg_1_43), .right(vreg_3_43), .up(vreg_2_44), .down(vreg_2_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_43), .sw(sw));
	wire signed[17:0] vwire_2_44;
	reg signed[17:0] vreg_2_44;
	node n2_44(.left(vreg_1_44), .right(vreg_3_44), .up(vreg_2_45), .down(vreg_2_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_44), .sw(sw));
	wire signed[17:0] vwire_2_45;
	reg signed[17:0] vreg_2_45;
	node n2_45(.left(vreg_1_45), .right(vreg_3_45), .up(vreg_2_46), .down(vreg_2_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_45), .sw(sw));
	wire signed[17:0] vwire_2_46;
	reg signed[17:0] vreg_2_46;
	node n2_46(.left(vreg_1_46), .right(vreg_3_46), .up(vreg_2_47), .down(vreg_2_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_46), .sw(sw));
	wire signed[17:0] vwire_2_47;
	reg signed[17:0] vreg_2_47;
	node n2_47(.left(vreg_1_47), .right(vreg_3_47), .up(vreg_2_48), .down(vreg_2_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_47), .sw(sw));
	wire signed[17:0] vwire_2_48;
	reg signed[17:0] vreg_2_48;
	node n2_48(.left(vreg_1_48), .right(vreg_3_48), .up(vreg_2_49), .down(vreg_2_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_48), .sw(sw));
	wire signed[17:0] vwire_2_49;
	reg signed[17:0] vreg_2_49;
	node n2_49(.left(vreg_1_49), .right(vreg_3_49), .up(18'b0), .down(vreg_2_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_49), .sw(sw));
	wire signed[17:0] vwire_3_0;
	reg signed[17:0] vreg_3_0;
	node n3_0(.left(vreg_2_0), .right(vreg_4_0), .up(vreg_3_1), .down(vreg_3_1), .clk(clk), .reset(restart), .resetval(18'b000000000111001111), .value(vwire_3_0), .sw(sw));
	wire signed[17:0] vwire_3_1;
	reg signed[17:0] vreg_3_1;
	node n3_1(.left(vreg_2_1), .right(vreg_4_1), .up(vreg_3_2), .down(vreg_3_0), .clk(clk), .reset(restart), .resetval(18'b000000000100011001), .value(vwire_3_1), .sw(sw));
	wire signed[17:0] vwire_3_2;
	reg signed[17:0] vreg_3_2;
	node n3_2(.left(vreg_2_2), .right(vreg_4_2), .up(vreg_3_3), .down(vreg_3_1), .clk(clk), .reset(restart), .resetval(18'b000000000000111111), .value(vwire_3_2), .sw(sw));
	wire signed[17:0] vwire_3_3;
	reg signed[17:0] vreg_3_3;
	node n3_3(.left(vreg_2_3), .right(vreg_4_3), .up(vreg_3_4), .down(vreg_3_2), .clk(clk), .reset(restart), .resetval(18'b000000000000000000), .value(vwire_3_3), .sw(sw));
	wire signed[17:0] vwire_3_4;
	reg signed[17:0] vreg_3_4;
	node n3_4(.left(vreg_2_4), .right(vreg_4_4), .up(vreg_3_5), .down(vreg_3_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_4), .sw(sw));
	wire signed[17:0] vwire_3_5;
	reg signed[17:0] vreg_3_5;
	node n3_5(.left(vreg_2_5), .right(vreg_4_5), .up(vreg_3_6), .down(vreg_3_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_5), .sw(sw));
	wire signed[17:0] vwire_3_6;
	reg signed[17:0] vreg_3_6;
	node n3_6(.left(vreg_2_6), .right(vreg_4_6), .up(vreg_3_7), .down(vreg_3_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_6), .sw(sw));
	wire signed[17:0] vwire_3_7;
	reg signed[17:0] vreg_3_7;
	node n3_7(.left(vreg_2_7), .right(vreg_4_7), .up(vreg_3_8), .down(vreg_3_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_7), .sw(sw));
	wire signed[17:0] vwire_3_8;
	reg signed[17:0] vreg_3_8;
	node n3_8(.left(vreg_2_8), .right(vreg_4_8), .up(vreg_3_9), .down(vreg_3_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_8), .sw(sw));
	wire signed[17:0] vwire_3_9;
	reg signed[17:0] vreg_3_9;
	node n3_9(.left(vreg_2_9), .right(vreg_4_9), .up(vreg_3_10), .down(vreg_3_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_9), .sw(sw));
	wire signed[17:0] vwire_3_10;
	reg signed[17:0] vreg_3_10;
	node n3_10(.left(vreg_2_10), .right(vreg_4_10), .up(vreg_3_11), .down(vreg_3_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_10), .sw(sw));
	wire signed[17:0] vwire_3_11;
	reg signed[17:0] vreg_3_11;
	node n3_11(.left(vreg_2_11), .right(vreg_4_11), .up(vreg_3_12), .down(vreg_3_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_11), .sw(sw));
	wire signed[17:0] vwire_3_12;
	reg signed[17:0] vreg_3_12;
	node n3_12(.left(vreg_2_12), .right(vreg_4_12), .up(vreg_3_13), .down(vreg_3_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_12), .sw(sw));
	wire signed[17:0] vwire_3_13;
	reg signed[17:0] vreg_3_13;
	node n3_13(.left(vreg_2_13), .right(vreg_4_13), .up(vreg_3_14), .down(vreg_3_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_13), .sw(sw));
	wire signed[17:0] vwire_3_14;
	reg signed[17:0] vreg_3_14;
	node n3_14(.left(vreg_2_14), .right(vreg_4_14), .up(vreg_3_15), .down(vreg_3_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_14), .sw(sw));
	wire signed[17:0] vwire_3_15;
	reg signed[17:0] vreg_3_15;
	node n3_15(.left(vreg_2_15), .right(vreg_4_15), .up(vreg_3_16), .down(vreg_3_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_15), .sw(sw));
	wire signed[17:0] vwire_3_16;
	reg signed[17:0] vreg_3_16;
	node n3_16(.left(vreg_2_16), .right(vreg_4_16), .up(vreg_3_17), .down(vreg_3_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_16), .sw(sw));
	wire signed[17:0] vwire_3_17;
	reg signed[17:0] vreg_3_17;
	node n3_17(.left(vreg_2_17), .right(vreg_4_17), .up(vreg_3_18), .down(vreg_3_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_17), .sw(sw));
	wire signed[17:0] vwire_3_18;
	reg signed[17:0] vreg_3_18;
	node n3_18(.left(vreg_2_18), .right(vreg_4_18), .up(vreg_3_19), .down(vreg_3_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_18), .sw(sw));
	wire signed[17:0] vwire_3_19;
	reg signed[17:0] vreg_3_19;
	node n3_19(.left(vreg_2_19), .right(vreg_4_19), .up(vreg_3_20), .down(vreg_3_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_19), .sw(sw));
	wire signed[17:0] vwire_3_20;
	reg signed[17:0] vreg_3_20;
	node n3_20(.left(vreg_2_20), .right(vreg_4_20), .up(vreg_3_21), .down(vreg_3_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_20), .sw(sw));
	wire signed[17:0] vwire_3_21;
	reg signed[17:0] vreg_3_21;
	node n3_21(.left(vreg_2_21), .right(vreg_4_21), .up(vreg_3_22), .down(vreg_3_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_21), .sw(sw));
	wire signed[17:0] vwire_3_22;
	reg signed[17:0] vreg_3_22;
	node n3_22(.left(vreg_2_22), .right(vreg_4_22), .up(vreg_3_23), .down(vreg_3_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_22), .sw(sw));
	wire signed[17:0] vwire_3_23;
	reg signed[17:0] vreg_3_23;
	node n3_23(.left(vreg_2_23), .right(vreg_4_23), .up(vreg_3_24), .down(vreg_3_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_23), .sw(sw));
	wire signed[17:0] vwire_3_24;
	reg signed[17:0] vreg_3_24;
	node n3_24(.left(vreg_2_24), .right(vreg_4_24), .up(vreg_3_25), .down(vreg_3_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_24), .sw(sw));
	wire signed[17:0] vwire_3_25;
	reg signed[17:0] vreg_3_25;
	node n3_25(.left(vreg_2_25), .right(vreg_4_25), .up(vreg_3_26), .down(vreg_3_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_25), .sw(sw));
	wire signed[17:0] vwire_3_26;
	reg signed[17:0] vreg_3_26;
	node n3_26(.left(vreg_2_26), .right(vreg_4_26), .up(vreg_3_27), .down(vreg_3_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_26), .sw(sw));
	wire signed[17:0] vwire_3_27;
	reg signed[17:0] vreg_3_27;
	node n3_27(.left(vreg_2_27), .right(vreg_4_27), .up(vreg_3_28), .down(vreg_3_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_27), .sw(sw));
	wire signed[17:0] vwire_3_28;
	reg signed[17:0] vreg_3_28;
	node n3_28(.left(vreg_2_28), .right(vreg_4_28), .up(vreg_3_29), .down(vreg_3_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_28), .sw(sw));
	wire signed[17:0] vwire_3_29;
	reg signed[17:0] vreg_3_29;
	node n3_29(.left(vreg_2_29), .right(vreg_4_29), .up(vreg_3_30), .down(vreg_3_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_29), .sw(sw));
	wire signed[17:0] vwire_3_30;
	reg signed[17:0] vreg_3_30;
	node n3_30(.left(vreg_2_30), .right(vreg_4_30), .up(vreg_3_31), .down(vreg_3_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_30), .sw(sw));
	wire signed[17:0] vwire_3_31;
	reg signed[17:0] vreg_3_31;
	node n3_31(.left(vreg_2_31), .right(vreg_4_31), .up(vreg_3_32), .down(vreg_3_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_31), .sw(sw));
	wire signed[17:0] vwire_3_32;
	reg signed[17:0] vreg_3_32;
	node n3_32(.left(vreg_2_32), .right(vreg_4_32), .up(vreg_3_33), .down(vreg_3_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_32), .sw(sw));
	wire signed[17:0] vwire_3_33;
	reg signed[17:0] vreg_3_33;
	node n3_33(.left(vreg_2_33), .right(vreg_4_33), .up(vreg_3_34), .down(vreg_3_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_33), .sw(sw));
	wire signed[17:0] vwire_3_34;
	reg signed[17:0] vreg_3_34;
	node n3_34(.left(vreg_2_34), .right(vreg_4_34), .up(vreg_3_35), .down(vreg_3_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_34), .sw(sw));
	wire signed[17:0] vwire_3_35;
	reg signed[17:0] vreg_3_35;
	node n3_35(.left(vreg_2_35), .right(vreg_4_35), .up(vreg_3_36), .down(vreg_3_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_35), .sw(sw));
	wire signed[17:0] vwire_3_36;
	reg signed[17:0] vreg_3_36;
	node n3_36(.left(vreg_2_36), .right(vreg_4_36), .up(vreg_3_37), .down(vreg_3_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_36), .sw(sw));
	wire signed[17:0] vwire_3_37;
	reg signed[17:0] vreg_3_37;
	node n3_37(.left(vreg_2_37), .right(vreg_4_37), .up(vreg_3_38), .down(vreg_3_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_37), .sw(sw));
	wire signed[17:0] vwire_3_38;
	reg signed[17:0] vreg_3_38;
	node n3_38(.left(vreg_2_38), .right(vreg_4_38), .up(vreg_3_39), .down(vreg_3_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_38), .sw(sw));
	wire signed[17:0] vwire_3_39;
	reg signed[17:0] vreg_3_39;
	node n3_39(.left(vreg_2_39), .right(vreg_4_39), .up(vreg_3_40), .down(vreg_3_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_39), .sw(sw));
	wire signed[17:0] vwire_3_40;
	reg signed[17:0] vreg_3_40;
	node n3_40(.left(vreg_2_40), .right(vreg_4_40), .up(vreg_3_41), .down(vreg_3_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_40), .sw(sw));
	wire signed[17:0] vwire_3_41;
	reg signed[17:0] vreg_3_41;
	node n3_41(.left(vreg_2_41), .right(vreg_4_41), .up(vreg_3_42), .down(vreg_3_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_41), .sw(sw));
	wire signed[17:0] vwire_3_42;
	reg signed[17:0] vreg_3_42;
	node n3_42(.left(vreg_2_42), .right(vreg_4_42), .up(vreg_3_43), .down(vreg_3_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_42), .sw(sw));
	wire signed[17:0] vwire_3_43;
	reg signed[17:0] vreg_3_43;
	node n3_43(.left(vreg_2_43), .right(vreg_4_43), .up(vreg_3_44), .down(vreg_3_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_43), .sw(sw));
	wire signed[17:0] vwire_3_44;
	reg signed[17:0] vreg_3_44;
	node n3_44(.left(vreg_2_44), .right(vreg_4_44), .up(vreg_3_45), .down(vreg_3_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_44), .sw(sw));
	wire signed[17:0] vwire_3_45;
	reg signed[17:0] vreg_3_45;
	node n3_45(.left(vreg_2_45), .right(vreg_4_45), .up(vreg_3_46), .down(vreg_3_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_45), .sw(sw));
	wire signed[17:0] vwire_3_46;
	reg signed[17:0] vreg_3_46;
	node n3_46(.left(vreg_2_46), .right(vreg_4_46), .up(vreg_3_47), .down(vreg_3_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_46), .sw(sw));
	wire signed[17:0] vwire_3_47;
	reg signed[17:0] vreg_3_47;
	node n3_47(.left(vreg_2_47), .right(vreg_4_47), .up(vreg_3_48), .down(vreg_3_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_47), .sw(sw));
	wire signed[17:0] vwire_3_48;
	reg signed[17:0] vreg_3_48;
	node n3_48(.left(vreg_2_48), .right(vreg_4_48), .up(vreg_3_49), .down(vreg_3_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_48), .sw(sw));
	wire signed[17:0] vwire_3_49;
	reg signed[17:0] vreg_3_49;
	node n3_49(.left(vreg_2_49), .right(vreg_4_49), .up(18'b0), .down(vreg_3_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_49), .sw(sw));
	wire signed[17:0] vwire_4_0;
	reg signed[17:0] vreg_4_0;
	node n4_0(.left(vreg_3_0), .right(vreg_5_0), .up(vreg_4_1), .down(vreg_4_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_0), .sw(sw));
	wire signed[17:0] vwire_4_1;
	reg signed[17:0] vreg_4_1;
	node n4_1(.left(vreg_3_1), .right(vreg_5_1), .up(vreg_4_2), .down(vreg_4_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_1), .sw(sw));
	wire signed[17:0] vwire_4_2;
	reg signed[17:0] vreg_4_2;
	node n4_2(.left(vreg_3_2), .right(vreg_5_2), .up(vreg_4_3), .down(vreg_4_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_2), .sw(sw));
	wire signed[17:0] vwire_4_3;
	reg signed[17:0] vreg_4_3;
	node n4_3(.left(vreg_3_3), .right(vreg_5_3), .up(vreg_4_4), .down(vreg_4_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_3), .sw(sw));
	wire signed[17:0] vwire_4_4;
	reg signed[17:0] vreg_4_4;
	node n4_4(.left(vreg_3_4), .right(vreg_5_4), .up(vreg_4_5), .down(vreg_4_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_4), .sw(sw));
	wire signed[17:0] vwire_4_5;
	reg signed[17:0] vreg_4_5;
	node n4_5(.left(vreg_3_5), .right(vreg_5_5), .up(vreg_4_6), .down(vreg_4_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_5), .sw(sw));
	wire signed[17:0] vwire_4_6;
	reg signed[17:0] vreg_4_6;
	node n4_6(.left(vreg_3_6), .right(vreg_5_6), .up(vreg_4_7), .down(vreg_4_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_6), .sw(sw));
	wire signed[17:0] vwire_4_7;
	reg signed[17:0] vreg_4_7;
	node n4_7(.left(vreg_3_7), .right(vreg_5_7), .up(vreg_4_8), .down(vreg_4_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_7), .sw(sw));
	wire signed[17:0] vwire_4_8;
	reg signed[17:0] vreg_4_8;
	node n4_8(.left(vreg_3_8), .right(vreg_5_8), .up(vreg_4_9), .down(vreg_4_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_8), .sw(sw));
	wire signed[17:0] vwire_4_9;
	reg signed[17:0] vreg_4_9;
	node n4_9(.left(vreg_3_9), .right(vreg_5_9), .up(vreg_4_10), .down(vreg_4_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_9), .sw(sw));
	wire signed[17:0] vwire_4_10;
	reg signed[17:0] vreg_4_10;
	node n4_10(.left(vreg_3_10), .right(vreg_5_10), .up(vreg_4_11), .down(vreg_4_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_10), .sw(sw));
	wire signed[17:0] vwire_4_11;
	reg signed[17:0] vreg_4_11;
	node n4_11(.left(vreg_3_11), .right(vreg_5_11), .up(vreg_4_12), .down(vreg_4_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_11), .sw(sw));
	wire signed[17:0] vwire_4_12;
	reg signed[17:0] vreg_4_12;
	node n4_12(.left(vreg_3_12), .right(vreg_5_12), .up(vreg_4_13), .down(vreg_4_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_12), .sw(sw));
	wire signed[17:0] vwire_4_13;
	reg signed[17:0] vreg_4_13;
	node n4_13(.left(vreg_3_13), .right(vreg_5_13), .up(vreg_4_14), .down(vreg_4_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_13), .sw(sw));
	wire signed[17:0] vwire_4_14;
	reg signed[17:0] vreg_4_14;
	node n4_14(.left(vreg_3_14), .right(vreg_5_14), .up(vreg_4_15), .down(vreg_4_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_14), .sw(sw));
	wire signed[17:0] vwire_4_15;
	reg signed[17:0] vreg_4_15;
	node n4_15(.left(vreg_3_15), .right(vreg_5_15), .up(vreg_4_16), .down(vreg_4_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_15), .sw(sw));
	wire signed[17:0] vwire_4_16;
	reg signed[17:0] vreg_4_16;
	node n4_16(.left(vreg_3_16), .right(vreg_5_16), .up(vreg_4_17), .down(vreg_4_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_16), .sw(sw));
	wire signed[17:0] vwire_4_17;
	reg signed[17:0] vreg_4_17;
	node n4_17(.left(vreg_3_17), .right(vreg_5_17), .up(vreg_4_18), .down(vreg_4_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_17), .sw(sw));
	wire signed[17:0] vwire_4_18;
	reg signed[17:0] vreg_4_18;
	node n4_18(.left(vreg_3_18), .right(vreg_5_18), .up(vreg_4_19), .down(vreg_4_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_18), .sw(sw));
	wire signed[17:0] vwire_4_19;
	reg signed[17:0] vreg_4_19;
	node n4_19(.left(vreg_3_19), .right(vreg_5_19), .up(vreg_4_20), .down(vreg_4_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_19), .sw(sw));
	wire signed[17:0] vwire_4_20;
	reg signed[17:0] vreg_4_20;
	node n4_20(.left(vreg_3_20), .right(vreg_5_20), .up(vreg_4_21), .down(vreg_4_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_20), .sw(sw));
	wire signed[17:0] vwire_4_21;
	reg signed[17:0] vreg_4_21;
	node n4_21(.left(vreg_3_21), .right(vreg_5_21), .up(vreg_4_22), .down(vreg_4_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_21), .sw(sw));
	wire signed[17:0] vwire_4_22;
	reg signed[17:0] vreg_4_22;
	node n4_22(.left(vreg_3_22), .right(vreg_5_22), .up(vreg_4_23), .down(vreg_4_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_22), .sw(sw));
	wire signed[17:0] vwire_4_23;
	reg signed[17:0] vreg_4_23;
	node n4_23(.left(vreg_3_23), .right(vreg_5_23), .up(vreg_4_24), .down(vreg_4_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_23), .sw(sw));
	wire signed[17:0] vwire_4_24;
	reg signed[17:0] vreg_4_24;
	node n4_24(.left(vreg_3_24), .right(vreg_5_24), .up(vreg_4_25), .down(vreg_4_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_24), .sw(sw));
	wire signed[17:0] vwire_4_25;
	reg signed[17:0] vreg_4_25;
	node n4_25(.left(vreg_3_25), .right(vreg_5_25), .up(vreg_4_26), .down(vreg_4_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_25), .sw(sw));
	wire signed[17:0] vwire_4_26;
	reg signed[17:0] vreg_4_26;
	node n4_26(.left(vreg_3_26), .right(vreg_5_26), .up(vreg_4_27), .down(vreg_4_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_26), .sw(sw));
	wire signed[17:0] vwire_4_27;
	reg signed[17:0] vreg_4_27;
	node n4_27(.left(vreg_3_27), .right(vreg_5_27), .up(vreg_4_28), .down(vreg_4_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_27), .sw(sw));
	wire signed[17:0] vwire_4_28;
	reg signed[17:0] vreg_4_28;
	node n4_28(.left(vreg_3_28), .right(vreg_5_28), .up(vreg_4_29), .down(vreg_4_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_28), .sw(sw));
	wire signed[17:0] vwire_4_29;
	reg signed[17:0] vreg_4_29;
	node n4_29(.left(vreg_3_29), .right(vreg_5_29), .up(vreg_4_30), .down(vreg_4_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_29), .sw(sw));
	wire signed[17:0] vwire_4_30;
	reg signed[17:0] vreg_4_30;
	node n4_30(.left(vreg_3_30), .right(vreg_5_30), .up(vreg_4_31), .down(vreg_4_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_30), .sw(sw));
	wire signed[17:0] vwire_4_31;
	reg signed[17:0] vreg_4_31;
	node n4_31(.left(vreg_3_31), .right(vreg_5_31), .up(vreg_4_32), .down(vreg_4_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_31), .sw(sw));
	wire signed[17:0] vwire_4_32;
	reg signed[17:0] vreg_4_32;
	node n4_32(.left(vreg_3_32), .right(vreg_5_32), .up(vreg_4_33), .down(vreg_4_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_32), .sw(sw));
	wire signed[17:0] vwire_4_33;
	reg signed[17:0] vreg_4_33;
	node n4_33(.left(vreg_3_33), .right(vreg_5_33), .up(vreg_4_34), .down(vreg_4_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_33), .sw(sw));
	wire signed[17:0] vwire_4_34;
	reg signed[17:0] vreg_4_34;
	node n4_34(.left(vreg_3_34), .right(vreg_5_34), .up(vreg_4_35), .down(vreg_4_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_34), .sw(sw));
	wire signed[17:0] vwire_4_35;
	reg signed[17:0] vreg_4_35;
	node n4_35(.left(vreg_3_35), .right(vreg_5_35), .up(vreg_4_36), .down(vreg_4_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_35), .sw(sw));
	wire signed[17:0] vwire_4_36;
	reg signed[17:0] vreg_4_36;
	node n4_36(.left(vreg_3_36), .right(vreg_5_36), .up(vreg_4_37), .down(vreg_4_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_36), .sw(sw));
	wire signed[17:0] vwire_4_37;
	reg signed[17:0] vreg_4_37;
	node n4_37(.left(vreg_3_37), .right(vreg_5_37), .up(vreg_4_38), .down(vreg_4_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_37), .sw(sw));
	wire signed[17:0] vwire_4_38;
	reg signed[17:0] vreg_4_38;
	node n4_38(.left(vreg_3_38), .right(vreg_5_38), .up(vreg_4_39), .down(vreg_4_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_38), .sw(sw));
	wire signed[17:0] vwire_4_39;
	reg signed[17:0] vreg_4_39;
	node n4_39(.left(vreg_3_39), .right(vreg_5_39), .up(vreg_4_40), .down(vreg_4_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_39), .sw(sw));
	wire signed[17:0] vwire_4_40;
	reg signed[17:0] vreg_4_40;
	node n4_40(.left(vreg_3_40), .right(vreg_5_40), .up(vreg_4_41), .down(vreg_4_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_40), .sw(sw));
	wire signed[17:0] vwire_4_41;
	reg signed[17:0] vreg_4_41;
	node n4_41(.left(vreg_3_41), .right(vreg_5_41), .up(vreg_4_42), .down(vreg_4_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_41), .sw(sw));
	wire signed[17:0] vwire_4_42;
	reg signed[17:0] vreg_4_42;
	node n4_42(.left(vreg_3_42), .right(vreg_5_42), .up(vreg_4_43), .down(vreg_4_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_42), .sw(sw));
	wire signed[17:0] vwire_4_43;
	reg signed[17:0] vreg_4_43;
	node n4_43(.left(vreg_3_43), .right(vreg_5_43), .up(vreg_4_44), .down(vreg_4_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_43), .sw(sw));
	wire signed[17:0] vwire_4_44;
	reg signed[17:0] vreg_4_44;
	node n4_44(.left(vreg_3_44), .right(vreg_5_44), .up(vreg_4_45), .down(vreg_4_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_44), .sw(sw));
	wire signed[17:0] vwire_4_45;
	reg signed[17:0] vreg_4_45;
	node n4_45(.left(vreg_3_45), .right(vreg_5_45), .up(vreg_4_46), .down(vreg_4_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_45), .sw(sw));
	wire signed[17:0] vwire_4_46;
	reg signed[17:0] vreg_4_46;
	node n4_46(.left(vreg_3_46), .right(vreg_5_46), .up(vreg_4_47), .down(vreg_4_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_46), .sw(sw));
	wire signed[17:0] vwire_4_47;
	reg signed[17:0] vreg_4_47;
	node n4_47(.left(vreg_3_47), .right(vreg_5_47), .up(vreg_4_48), .down(vreg_4_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_47), .sw(sw));
	wire signed[17:0] vwire_4_48;
	reg signed[17:0] vreg_4_48;
	node n4_48(.left(vreg_3_48), .right(vreg_5_48), .up(vreg_4_49), .down(vreg_4_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_48), .sw(sw));
	wire signed[17:0] vwire_4_49;
	reg signed[17:0] vreg_4_49;
	node n4_49(.left(vreg_3_49), .right(vreg_5_49), .up(18'b0), .down(vreg_4_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_49), .sw(sw));
	wire signed[17:0] vwire_5_0;
	reg signed[17:0] vreg_5_0;
	node n5_0(.left(vreg_4_0), .right(vreg_6_0), .up(vreg_5_1), .down(vreg_5_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_0), .sw(sw));
	wire signed[17:0] vwire_5_1;
	reg signed[17:0] vreg_5_1;
	node n5_1(.left(vreg_4_1), .right(vreg_6_1), .up(vreg_5_2), .down(vreg_5_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_1), .sw(sw));
	wire signed[17:0] vwire_5_2;
	reg signed[17:0] vreg_5_2;
	node n5_2(.left(vreg_4_2), .right(vreg_6_2), .up(vreg_5_3), .down(vreg_5_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_2), .sw(sw));
	wire signed[17:0] vwire_5_3;
	reg signed[17:0] vreg_5_3;
	node n5_3(.left(vreg_4_3), .right(vreg_6_3), .up(vreg_5_4), .down(vreg_5_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_3), .sw(sw));
	wire signed[17:0] vwire_5_4;
	reg signed[17:0] vreg_5_4;
	node n5_4(.left(vreg_4_4), .right(vreg_6_4), .up(vreg_5_5), .down(vreg_5_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_4), .sw(sw));
	wire signed[17:0] vwire_5_5;
	reg signed[17:0] vreg_5_5;
	node n5_5(.left(vreg_4_5), .right(vreg_6_5), .up(vreg_5_6), .down(vreg_5_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_5), .sw(sw));
	wire signed[17:0] vwire_5_6;
	reg signed[17:0] vreg_5_6;
	node n5_6(.left(vreg_4_6), .right(vreg_6_6), .up(vreg_5_7), .down(vreg_5_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_6), .sw(sw));
	wire signed[17:0] vwire_5_7;
	reg signed[17:0] vreg_5_7;
	node n5_7(.left(vreg_4_7), .right(vreg_6_7), .up(vreg_5_8), .down(vreg_5_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_7), .sw(sw));
	wire signed[17:0] vwire_5_8;
	reg signed[17:0] vreg_5_8;
	node n5_8(.left(vreg_4_8), .right(vreg_6_8), .up(vreg_5_9), .down(vreg_5_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_8), .sw(sw));
	wire signed[17:0] vwire_5_9;
	reg signed[17:0] vreg_5_9;
	node n5_9(.left(vreg_4_9), .right(vreg_6_9), .up(vreg_5_10), .down(vreg_5_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_9), .sw(sw));
	wire signed[17:0] vwire_5_10;
	reg signed[17:0] vreg_5_10;
	node n5_10(.left(vreg_4_10), .right(vreg_6_10), .up(vreg_5_11), .down(vreg_5_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_10), .sw(sw));
	wire signed[17:0] vwire_5_11;
	reg signed[17:0] vreg_5_11;
	node n5_11(.left(vreg_4_11), .right(vreg_6_11), .up(vreg_5_12), .down(vreg_5_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_11), .sw(sw));
	wire signed[17:0] vwire_5_12;
	reg signed[17:0] vreg_5_12;
	node n5_12(.left(vreg_4_12), .right(vreg_6_12), .up(vreg_5_13), .down(vreg_5_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_12), .sw(sw));
	wire signed[17:0] vwire_5_13;
	reg signed[17:0] vreg_5_13;
	node n5_13(.left(vreg_4_13), .right(vreg_6_13), .up(vreg_5_14), .down(vreg_5_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_13), .sw(sw));
	wire signed[17:0] vwire_5_14;
	reg signed[17:0] vreg_5_14;
	node n5_14(.left(vreg_4_14), .right(vreg_6_14), .up(vreg_5_15), .down(vreg_5_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_14), .sw(sw));
	wire signed[17:0] vwire_5_15;
	reg signed[17:0] vreg_5_15;
	node n5_15(.left(vreg_4_15), .right(vreg_6_15), .up(vreg_5_16), .down(vreg_5_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_15), .sw(sw));
	wire signed[17:0] vwire_5_16;
	reg signed[17:0] vreg_5_16;
	node n5_16(.left(vreg_4_16), .right(vreg_6_16), .up(vreg_5_17), .down(vreg_5_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_16), .sw(sw));
	wire signed[17:0] vwire_5_17;
	reg signed[17:0] vreg_5_17;
	node n5_17(.left(vreg_4_17), .right(vreg_6_17), .up(vreg_5_18), .down(vreg_5_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_17), .sw(sw));
	wire signed[17:0] vwire_5_18;
	reg signed[17:0] vreg_5_18;
	node n5_18(.left(vreg_4_18), .right(vreg_6_18), .up(vreg_5_19), .down(vreg_5_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_18), .sw(sw));
	wire signed[17:0] vwire_5_19;
	reg signed[17:0] vreg_5_19;
	node n5_19(.left(vreg_4_19), .right(vreg_6_19), .up(vreg_5_20), .down(vreg_5_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_19), .sw(sw));
	wire signed[17:0] vwire_5_20;
	reg signed[17:0] vreg_5_20;
	node n5_20(.left(vreg_4_20), .right(vreg_6_20), .up(vreg_5_21), .down(vreg_5_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_20), .sw(sw));
	wire signed[17:0] vwire_5_21;
	reg signed[17:0] vreg_5_21;
	node n5_21(.left(vreg_4_21), .right(vreg_6_21), .up(vreg_5_22), .down(vreg_5_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_21), .sw(sw));
	wire signed[17:0] vwire_5_22;
	reg signed[17:0] vreg_5_22;
	node n5_22(.left(vreg_4_22), .right(vreg_6_22), .up(vreg_5_23), .down(vreg_5_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_22), .sw(sw));
	wire signed[17:0] vwire_5_23;
	reg signed[17:0] vreg_5_23;
	node n5_23(.left(vreg_4_23), .right(vreg_6_23), .up(vreg_5_24), .down(vreg_5_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_23), .sw(sw));
	wire signed[17:0] vwire_5_24;
	reg signed[17:0] vreg_5_24;
	node n5_24(.left(vreg_4_24), .right(vreg_6_24), .up(vreg_5_25), .down(vreg_5_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_24), .sw(sw));
	wire signed[17:0] vwire_5_25;
	reg signed[17:0] vreg_5_25;
	node n5_25(.left(vreg_4_25), .right(vreg_6_25), .up(vreg_5_26), .down(vreg_5_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_25), .sw(sw));
	wire signed[17:0] vwire_5_26;
	reg signed[17:0] vreg_5_26;
	node n5_26(.left(vreg_4_26), .right(vreg_6_26), .up(vreg_5_27), .down(vreg_5_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_26), .sw(sw));
	wire signed[17:0] vwire_5_27;
	reg signed[17:0] vreg_5_27;
	node n5_27(.left(vreg_4_27), .right(vreg_6_27), .up(vreg_5_28), .down(vreg_5_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_27), .sw(sw));
	wire signed[17:0] vwire_5_28;
	reg signed[17:0] vreg_5_28;
	node n5_28(.left(vreg_4_28), .right(vreg_6_28), .up(vreg_5_29), .down(vreg_5_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_28), .sw(sw));
	wire signed[17:0] vwire_5_29;
	reg signed[17:0] vreg_5_29;
	node n5_29(.left(vreg_4_29), .right(vreg_6_29), .up(vreg_5_30), .down(vreg_5_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_29), .sw(sw));
	wire signed[17:0] vwire_5_30;
	reg signed[17:0] vreg_5_30;
	node n5_30(.left(vreg_4_30), .right(vreg_6_30), .up(vreg_5_31), .down(vreg_5_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_30), .sw(sw));
	wire signed[17:0] vwire_5_31;
	reg signed[17:0] vreg_5_31;
	node n5_31(.left(vreg_4_31), .right(vreg_6_31), .up(vreg_5_32), .down(vreg_5_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_31), .sw(sw));
	wire signed[17:0] vwire_5_32;
	reg signed[17:0] vreg_5_32;
	node n5_32(.left(vreg_4_32), .right(vreg_6_32), .up(vreg_5_33), .down(vreg_5_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_32), .sw(sw));
	wire signed[17:0] vwire_5_33;
	reg signed[17:0] vreg_5_33;
	node n5_33(.left(vreg_4_33), .right(vreg_6_33), .up(vreg_5_34), .down(vreg_5_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_33), .sw(sw));
	wire signed[17:0] vwire_5_34;
	reg signed[17:0] vreg_5_34;
	node n5_34(.left(vreg_4_34), .right(vreg_6_34), .up(vreg_5_35), .down(vreg_5_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_34), .sw(sw));
	wire signed[17:0] vwire_5_35;
	reg signed[17:0] vreg_5_35;
	node n5_35(.left(vreg_4_35), .right(vreg_6_35), .up(vreg_5_36), .down(vreg_5_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_35), .sw(sw));
	wire signed[17:0] vwire_5_36;
	reg signed[17:0] vreg_5_36;
	node n5_36(.left(vreg_4_36), .right(vreg_6_36), .up(vreg_5_37), .down(vreg_5_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_36), .sw(sw));
	wire signed[17:0] vwire_5_37;
	reg signed[17:0] vreg_5_37;
	node n5_37(.left(vreg_4_37), .right(vreg_6_37), .up(vreg_5_38), .down(vreg_5_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_37), .sw(sw));
	wire signed[17:0] vwire_5_38;
	reg signed[17:0] vreg_5_38;
	node n5_38(.left(vreg_4_38), .right(vreg_6_38), .up(vreg_5_39), .down(vreg_5_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_38), .sw(sw));
	wire signed[17:0] vwire_5_39;
	reg signed[17:0] vreg_5_39;
	node n5_39(.left(vreg_4_39), .right(vreg_6_39), .up(vreg_5_40), .down(vreg_5_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_39), .sw(sw));
	wire signed[17:0] vwire_5_40;
	reg signed[17:0] vreg_5_40;
	node n5_40(.left(vreg_4_40), .right(vreg_6_40), .up(vreg_5_41), .down(vreg_5_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_40), .sw(sw));
	wire signed[17:0] vwire_5_41;
	reg signed[17:0] vreg_5_41;
	node n5_41(.left(vreg_4_41), .right(vreg_6_41), .up(vreg_5_42), .down(vreg_5_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_41), .sw(sw));
	wire signed[17:0] vwire_5_42;
	reg signed[17:0] vreg_5_42;
	node n5_42(.left(vreg_4_42), .right(vreg_6_42), .up(vreg_5_43), .down(vreg_5_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_42), .sw(sw));
	wire signed[17:0] vwire_5_43;
	reg signed[17:0] vreg_5_43;
	node n5_43(.left(vreg_4_43), .right(vreg_6_43), .up(vreg_5_44), .down(vreg_5_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_43), .sw(sw));
	wire signed[17:0] vwire_5_44;
	reg signed[17:0] vreg_5_44;
	node n5_44(.left(vreg_4_44), .right(vreg_6_44), .up(vreg_5_45), .down(vreg_5_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_44), .sw(sw));
	wire signed[17:0] vwire_5_45;
	reg signed[17:0] vreg_5_45;
	node n5_45(.left(vreg_4_45), .right(vreg_6_45), .up(vreg_5_46), .down(vreg_5_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_45), .sw(sw));
	wire signed[17:0] vwire_5_46;
	reg signed[17:0] vreg_5_46;
	node n5_46(.left(vreg_4_46), .right(vreg_6_46), .up(vreg_5_47), .down(vreg_5_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_46), .sw(sw));
	wire signed[17:0] vwire_5_47;
	reg signed[17:0] vreg_5_47;
	node n5_47(.left(vreg_4_47), .right(vreg_6_47), .up(vreg_5_48), .down(vreg_5_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_47), .sw(sw));
	wire signed[17:0] vwire_5_48;
	reg signed[17:0] vreg_5_48;
	node n5_48(.left(vreg_4_48), .right(vreg_6_48), .up(vreg_5_49), .down(vreg_5_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_48), .sw(sw));
	wire signed[17:0] vwire_5_49;
	reg signed[17:0] vreg_5_49;
	node n5_49(.left(vreg_4_49), .right(vreg_6_49), .up(18'b0), .down(vreg_5_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_49), .sw(sw));
	wire signed[17:0] vwire_6_0;
	reg signed[17:0] vreg_6_0;
	node n6_0(.left(vreg_5_0), .right(vreg_7_0), .up(vreg_6_1), .down(vreg_6_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_0), .sw(sw));
	wire signed[17:0] vwire_6_1;
	reg signed[17:0] vreg_6_1;
	node n6_1(.left(vreg_5_1), .right(vreg_7_1), .up(vreg_6_2), .down(vreg_6_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_1), .sw(sw));
	wire signed[17:0] vwire_6_2;
	reg signed[17:0] vreg_6_2;
	node n6_2(.left(vreg_5_2), .right(vreg_7_2), .up(vreg_6_3), .down(vreg_6_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_2), .sw(sw));
	wire signed[17:0] vwire_6_3;
	reg signed[17:0] vreg_6_3;
	node n6_3(.left(vreg_5_3), .right(vreg_7_3), .up(vreg_6_4), .down(vreg_6_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_3), .sw(sw));
	wire signed[17:0] vwire_6_4;
	reg signed[17:0] vreg_6_4;
	node n6_4(.left(vreg_5_4), .right(vreg_7_4), .up(vreg_6_5), .down(vreg_6_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_4), .sw(sw));
	wire signed[17:0] vwire_6_5;
	reg signed[17:0] vreg_6_5;
	node n6_5(.left(vreg_5_5), .right(vreg_7_5), .up(vreg_6_6), .down(vreg_6_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_5), .sw(sw));
	wire signed[17:0] vwire_6_6;
	reg signed[17:0] vreg_6_6;
	node n6_6(.left(vreg_5_6), .right(vreg_7_6), .up(vreg_6_7), .down(vreg_6_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_6), .sw(sw));
	wire signed[17:0] vwire_6_7;
	reg signed[17:0] vreg_6_7;
	node n6_7(.left(vreg_5_7), .right(vreg_7_7), .up(vreg_6_8), .down(vreg_6_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_7), .sw(sw));
	wire signed[17:0] vwire_6_8;
	reg signed[17:0] vreg_6_8;
	node n6_8(.left(vreg_5_8), .right(vreg_7_8), .up(vreg_6_9), .down(vreg_6_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_8), .sw(sw));
	wire signed[17:0] vwire_6_9;
	reg signed[17:0] vreg_6_9;
	node n6_9(.left(vreg_5_9), .right(vreg_7_9), .up(vreg_6_10), .down(vreg_6_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_9), .sw(sw));
	wire signed[17:0] vwire_6_10;
	reg signed[17:0] vreg_6_10;
	node n6_10(.left(vreg_5_10), .right(vreg_7_10), .up(vreg_6_11), .down(vreg_6_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_10), .sw(sw));
	wire signed[17:0] vwire_6_11;
	reg signed[17:0] vreg_6_11;
	node n6_11(.left(vreg_5_11), .right(vreg_7_11), .up(vreg_6_12), .down(vreg_6_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_11), .sw(sw));
	wire signed[17:0] vwire_6_12;
	reg signed[17:0] vreg_6_12;
	node n6_12(.left(vreg_5_12), .right(vreg_7_12), .up(vreg_6_13), .down(vreg_6_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_12), .sw(sw));
	wire signed[17:0] vwire_6_13;
	reg signed[17:0] vreg_6_13;
	node n6_13(.left(vreg_5_13), .right(vreg_7_13), .up(vreg_6_14), .down(vreg_6_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_13), .sw(sw));
	wire signed[17:0] vwire_6_14;
	reg signed[17:0] vreg_6_14;
	node n6_14(.left(vreg_5_14), .right(vreg_7_14), .up(vreg_6_15), .down(vreg_6_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_14), .sw(sw));
	wire signed[17:0] vwire_6_15;
	reg signed[17:0] vreg_6_15;
	node n6_15(.left(vreg_5_15), .right(vreg_7_15), .up(vreg_6_16), .down(vreg_6_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_15), .sw(sw));
	wire signed[17:0] vwire_6_16;
	reg signed[17:0] vreg_6_16;
	node n6_16(.left(vreg_5_16), .right(vreg_7_16), .up(vreg_6_17), .down(vreg_6_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_16), .sw(sw));
	wire signed[17:0] vwire_6_17;
	reg signed[17:0] vreg_6_17;
	node n6_17(.left(vreg_5_17), .right(vreg_7_17), .up(vreg_6_18), .down(vreg_6_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_17), .sw(sw));
	wire signed[17:0] vwire_6_18;
	reg signed[17:0] vreg_6_18;
	node n6_18(.left(vreg_5_18), .right(vreg_7_18), .up(vreg_6_19), .down(vreg_6_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_18), .sw(sw));
	wire signed[17:0] vwire_6_19;
	reg signed[17:0] vreg_6_19;
	node n6_19(.left(vreg_5_19), .right(vreg_7_19), .up(vreg_6_20), .down(vreg_6_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_19), .sw(sw));
	wire signed[17:0] vwire_6_20;
	reg signed[17:0] vreg_6_20;
	node n6_20(.left(vreg_5_20), .right(vreg_7_20), .up(vreg_6_21), .down(vreg_6_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_20), .sw(sw));
	wire signed[17:0] vwire_6_21;
	reg signed[17:0] vreg_6_21;
	node n6_21(.left(vreg_5_21), .right(vreg_7_21), .up(vreg_6_22), .down(vreg_6_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_21), .sw(sw));
	wire signed[17:0] vwire_6_22;
	reg signed[17:0] vreg_6_22;
	node n6_22(.left(vreg_5_22), .right(vreg_7_22), .up(vreg_6_23), .down(vreg_6_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_22), .sw(sw));
	wire signed[17:0] vwire_6_23;
	reg signed[17:0] vreg_6_23;
	node n6_23(.left(vreg_5_23), .right(vreg_7_23), .up(vreg_6_24), .down(vreg_6_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_23), .sw(sw));
	wire signed[17:0] vwire_6_24;
	reg signed[17:0] vreg_6_24;
	node n6_24(.left(vreg_5_24), .right(vreg_7_24), .up(vreg_6_25), .down(vreg_6_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_24), .sw(sw));
	wire signed[17:0] vwire_6_25;
	reg signed[17:0] vreg_6_25;
	node n6_25(.left(vreg_5_25), .right(vreg_7_25), .up(vreg_6_26), .down(vreg_6_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_25), .sw(sw));
	wire signed[17:0] vwire_6_26;
	reg signed[17:0] vreg_6_26;
	node n6_26(.left(vreg_5_26), .right(vreg_7_26), .up(vreg_6_27), .down(vreg_6_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_26), .sw(sw));
	wire signed[17:0] vwire_6_27;
	reg signed[17:0] vreg_6_27;
	node n6_27(.left(vreg_5_27), .right(vreg_7_27), .up(vreg_6_28), .down(vreg_6_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_27), .sw(sw));
	wire signed[17:0] vwire_6_28;
	reg signed[17:0] vreg_6_28;
	node n6_28(.left(vreg_5_28), .right(vreg_7_28), .up(vreg_6_29), .down(vreg_6_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_28), .sw(sw));
	wire signed[17:0] vwire_6_29;
	reg signed[17:0] vreg_6_29;
	node n6_29(.left(vreg_5_29), .right(vreg_7_29), .up(vreg_6_30), .down(vreg_6_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_29), .sw(sw));
	wire signed[17:0] vwire_6_30;
	reg signed[17:0] vreg_6_30;
	node n6_30(.left(vreg_5_30), .right(vreg_7_30), .up(vreg_6_31), .down(vreg_6_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_30), .sw(sw));
	wire signed[17:0] vwire_6_31;
	reg signed[17:0] vreg_6_31;
	node n6_31(.left(vreg_5_31), .right(vreg_7_31), .up(vreg_6_32), .down(vreg_6_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_31), .sw(sw));
	wire signed[17:0] vwire_6_32;
	reg signed[17:0] vreg_6_32;
	node n6_32(.left(vreg_5_32), .right(vreg_7_32), .up(vreg_6_33), .down(vreg_6_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_32), .sw(sw));
	wire signed[17:0] vwire_6_33;
	reg signed[17:0] vreg_6_33;
	node n6_33(.left(vreg_5_33), .right(vreg_7_33), .up(vreg_6_34), .down(vreg_6_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_33), .sw(sw));
	wire signed[17:0] vwire_6_34;
	reg signed[17:0] vreg_6_34;
	node n6_34(.left(vreg_5_34), .right(vreg_7_34), .up(vreg_6_35), .down(vreg_6_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_34), .sw(sw));
	wire signed[17:0] vwire_6_35;
	reg signed[17:0] vreg_6_35;
	node n6_35(.left(vreg_5_35), .right(vreg_7_35), .up(vreg_6_36), .down(vreg_6_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_35), .sw(sw));
	wire signed[17:0] vwire_6_36;
	reg signed[17:0] vreg_6_36;
	node n6_36(.left(vreg_5_36), .right(vreg_7_36), .up(vreg_6_37), .down(vreg_6_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_36), .sw(sw));
	wire signed[17:0] vwire_6_37;
	reg signed[17:0] vreg_6_37;
	node n6_37(.left(vreg_5_37), .right(vreg_7_37), .up(vreg_6_38), .down(vreg_6_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_37), .sw(sw));
	wire signed[17:0] vwire_6_38;
	reg signed[17:0] vreg_6_38;
	node n6_38(.left(vreg_5_38), .right(vreg_7_38), .up(vreg_6_39), .down(vreg_6_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_38), .sw(sw));
	wire signed[17:0] vwire_6_39;
	reg signed[17:0] vreg_6_39;
	node n6_39(.left(vreg_5_39), .right(vreg_7_39), .up(vreg_6_40), .down(vreg_6_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_39), .sw(sw));
	wire signed[17:0] vwire_6_40;
	reg signed[17:0] vreg_6_40;
	node n6_40(.left(vreg_5_40), .right(vreg_7_40), .up(vreg_6_41), .down(vreg_6_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_40), .sw(sw));
	wire signed[17:0] vwire_6_41;
	reg signed[17:0] vreg_6_41;
	node n6_41(.left(vreg_5_41), .right(vreg_7_41), .up(vreg_6_42), .down(vreg_6_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_41), .sw(sw));
	wire signed[17:0] vwire_6_42;
	reg signed[17:0] vreg_6_42;
	node n6_42(.left(vreg_5_42), .right(vreg_7_42), .up(vreg_6_43), .down(vreg_6_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_42), .sw(sw));
	wire signed[17:0] vwire_6_43;
	reg signed[17:0] vreg_6_43;
	node n6_43(.left(vreg_5_43), .right(vreg_7_43), .up(vreg_6_44), .down(vreg_6_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_43), .sw(sw));
	wire signed[17:0] vwire_6_44;
	reg signed[17:0] vreg_6_44;
	node n6_44(.left(vreg_5_44), .right(vreg_7_44), .up(vreg_6_45), .down(vreg_6_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_44), .sw(sw));
	wire signed[17:0] vwire_6_45;
	reg signed[17:0] vreg_6_45;
	node n6_45(.left(vreg_5_45), .right(vreg_7_45), .up(vreg_6_46), .down(vreg_6_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_45), .sw(sw));
	wire signed[17:0] vwire_6_46;
	reg signed[17:0] vreg_6_46;
	node n6_46(.left(vreg_5_46), .right(vreg_7_46), .up(vreg_6_47), .down(vreg_6_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_46), .sw(sw));
	wire signed[17:0] vwire_6_47;
	reg signed[17:0] vreg_6_47;
	node n6_47(.left(vreg_5_47), .right(vreg_7_47), .up(vreg_6_48), .down(vreg_6_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_47), .sw(sw));
	wire signed[17:0] vwire_6_48;
	reg signed[17:0] vreg_6_48;
	node n6_48(.left(vreg_5_48), .right(vreg_7_48), .up(vreg_6_49), .down(vreg_6_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_48), .sw(sw));
	wire signed[17:0] vwire_6_49;
	reg signed[17:0] vreg_6_49;
	node n6_49(.left(vreg_5_49), .right(vreg_7_49), .up(18'b0), .down(vreg_6_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_49), .sw(sw));
	wire signed[17:0] vwire_7_0;
	reg signed[17:0] vreg_7_0;
	node n7_0(.left(vreg_6_0), .right(vreg_8_0), .up(vreg_7_1), .down(vreg_7_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_0), .sw(sw));
	wire signed[17:0] vwire_7_1;
	reg signed[17:0] vreg_7_1;
	node n7_1(.left(vreg_6_1), .right(vreg_8_1), .up(vreg_7_2), .down(vreg_7_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_1), .sw(sw));
	wire signed[17:0] vwire_7_2;
	reg signed[17:0] vreg_7_2;
	node n7_2(.left(vreg_6_2), .right(vreg_8_2), .up(vreg_7_3), .down(vreg_7_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_2), .sw(sw));
	wire signed[17:0] vwire_7_3;
	reg signed[17:0] vreg_7_3;
	node n7_3(.left(vreg_6_3), .right(vreg_8_3), .up(vreg_7_4), .down(vreg_7_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_3), .sw(sw));
	wire signed[17:0] vwire_7_4;
	reg signed[17:0] vreg_7_4;
	node n7_4(.left(vreg_6_4), .right(vreg_8_4), .up(vreg_7_5), .down(vreg_7_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_4), .sw(sw));
	wire signed[17:0] vwire_7_5;
	reg signed[17:0] vreg_7_5;
	node n7_5(.left(vreg_6_5), .right(vreg_8_5), .up(vreg_7_6), .down(vreg_7_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_5), .sw(sw));
	wire signed[17:0] vwire_7_6;
	reg signed[17:0] vreg_7_6;
	node n7_6(.left(vreg_6_6), .right(vreg_8_6), .up(vreg_7_7), .down(vreg_7_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_6), .sw(sw));
	wire signed[17:0] vwire_7_7;
	reg signed[17:0] vreg_7_7;
	node n7_7(.left(vreg_6_7), .right(vreg_8_7), .up(vreg_7_8), .down(vreg_7_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_7), .sw(sw));
	wire signed[17:0] vwire_7_8;
	reg signed[17:0] vreg_7_8;
	node n7_8(.left(vreg_6_8), .right(vreg_8_8), .up(vreg_7_9), .down(vreg_7_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_8), .sw(sw));
	wire signed[17:0] vwire_7_9;
	reg signed[17:0] vreg_7_9;
	node n7_9(.left(vreg_6_9), .right(vreg_8_9), .up(vreg_7_10), .down(vreg_7_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_9), .sw(sw));
	wire signed[17:0] vwire_7_10;
	reg signed[17:0] vreg_7_10;
	node n7_10(.left(vreg_6_10), .right(vreg_8_10), .up(vreg_7_11), .down(vreg_7_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_10), .sw(sw));
	wire signed[17:0] vwire_7_11;
	reg signed[17:0] vreg_7_11;
	node n7_11(.left(vreg_6_11), .right(vreg_8_11), .up(vreg_7_12), .down(vreg_7_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_11), .sw(sw));
	wire signed[17:0] vwire_7_12;
	reg signed[17:0] vreg_7_12;
	node n7_12(.left(vreg_6_12), .right(vreg_8_12), .up(vreg_7_13), .down(vreg_7_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_12), .sw(sw));
	wire signed[17:0] vwire_7_13;
	reg signed[17:0] vreg_7_13;
	node n7_13(.left(vreg_6_13), .right(vreg_8_13), .up(vreg_7_14), .down(vreg_7_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_13), .sw(sw));
	wire signed[17:0] vwire_7_14;
	reg signed[17:0] vreg_7_14;
	node n7_14(.left(vreg_6_14), .right(vreg_8_14), .up(vreg_7_15), .down(vreg_7_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_14), .sw(sw));
	wire signed[17:0] vwire_7_15;
	reg signed[17:0] vreg_7_15;
	node n7_15(.left(vreg_6_15), .right(vreg_8_15), .up(vreg_7_16), .down(vreg_7_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_15), .sw(sw));
	wire signed[17:0] vwire_7_16;
	reg signed[17:0] vreg_7_16;
	node n7_16(.left(vreg_6_16), .right(vreg_8_16), .up(vreg_7_17), .down(vreg_7_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_16), .sw(sw));
	wire signed[17:0] vwire_7_17;
	reg signed[17:0] vreg_7_17;
	node n7_17(.left(vreg_6_17), .right(vreg_8_17), .up(vreg_7_18), .down(vreg_7_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_17), .sw(sw));
	wire signed[17:0] vwire_7_18;
	reg signed[17:0] vreg_7_18;
	node n7_18(.left(vreg_6_18), .right(vreg_8_18), .up(vreg_7_19), .down(vreg_7_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_18), .sw(sw));
	wire signed[17:0] vwire_7_19;
	reg signed[17:0] vreg_7_19;
	node n7_19(.left(vreg_6_19), .right(vreg_8_19), .up(vreg_7_20), .down(vreg_7_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_19), .sw(sw));
	wire signed[17:0] vwire_7_20;
	reg signed[17:0] vreg_7_20;
	node n7_20(.left(vreg_6_20), .right(vreg_8_20), .up(vreg_7_21), .down(vreg_7_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_20), .sw(sw));
	wire signed[17:0] vwire_7_21;
	reg signed[17:0] vreg_7_21;
	node n7_21(.left(vreg_6_21), .right(vreg_8_21), .up(vreg_7_22), .down(vreg_7_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_21), .sw(sw));
	wire signed[17:0] vwire_7_22;
	reg signed[17:0] vreg_7_22;
	node n7_22(.left(vreg_6_22), .right(vreg_8_22), .up(vreg_7_23), .down(vreg_7_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_22), .sw(sw));
	wire signed[17:0] vwire_7_23;
	reg signed[17:0] vreg_7_23;
	node n7_23(.left(vreg_6_23), .right(vreg_8_23), .up(vreg_7_24), .down(vreg_7_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_23), .sw(sw));
	wire signed[17:0] vwire_7_24;
	reg signed[17:0] vreg_7_24;
	node n7_24(.left(vreg_6_24), .right(vreg_8_24), .up(vreg_7_25), .down(vreg_7_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_24), .sw(sw));
	wire signed[17:0] vwire_7_25;
	reg signed[17:0] vreg_7_25;
	node n7_25(.left(vreg_6_25), .right(vreg_8_25), .up(vreg_7_26), .down(vreg_7_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_25), .sw(sw));
	wire signed[17:0] vwire_7_26;
	reg signed[17:0] vreg_7_26;
	node n7_26(.left(vreg_6_26), .right(vreg_8_26), .up(vreg_7_27), .down(vreg_7_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_26), .sw(sw));
	wire signed[17:0] vwire_7_27;
	reg signed[17:0] vreg_7_27;
	node n7_27(.left(vreg_6_27), .right(vreg_8_27), .up(vreg_7_28), .down(vreg_7_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_27), .sw(sw));
	wire signed[17:0] vwire_7_28;
	reg signed[17:0] vreg_7_28;
	node n7_28(.left(vreg_6_28), .right(vreg_8_28), .up(vreg_7_29), .down(vreg_7_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_28), .sw(sw));
	wire signed[17:0] vwire_7_29;
	reg signed[17:0] vreg_7_29;
	node n7_29(.left(vreg_6_29), .right(vreg_8_29), .up(vreg_7_30), .down(vreg_7_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_29), .sw(sw));
	wire signed[17:0] vwire_7_30;
	reg signed[17:0] vreg_7_30;
	node n7_30(.left(vreg_6_30), .right(vreg_8_30), .up(vreg_7_31), .down(vreg_7_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_30), .sw(sw));
	wire signed[17:0] vwire_7_31;
	reg signed[17:0] vreg_7_31;
	node n7_31(.left(vreg_6_31), .right(vreg_8_31), .up(vreg_7_32), .down(vreg_7_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_31), .sw(sw));
	wire signed[17:0] vwire_7_32;
	reg signed[17:0] vreg_7_32;
	node n7_32(.left(vreg_6_32), .right(vreg_8_32), .up(vreg_7_33), .down(vreg_7_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_32), .sw(sw));
	wire signed[17:0] vwire_7_33;
	reg signed[17:0] vreg_7_33;
	node n7_33(.left(vreg_6_33), .right(vreg_8_33), .up(vreg_7_34), .down(vreg_7_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_33), .sw(sw));
	wire signed[17:0] vwire_7_34;
	reg signed[17:0] vreg_7_34;
	node n7_34(.left(vreg_6_34), .right(vreg_8_34), .up(vreg_7_35), .down(vreg_7_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_34), .sw(sw));
	wire signed[17:0] vwire_7_35;
	reg signed[17:0] vreg_7_35;
	node n7_35(.left(vreg_6_35), .right(vreg_8_35), .up(vreg_7_36), .down(vreg_7_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_35), .sw(sw));
	wire signed[17:0] vwire_7_36;
	reg signed[17:0] vreg_7_36;
	node n7_36(.left(vreg_6_36), .right(vreg_8_36), .up(vreg_7_37), .down(vreg_7_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_36), .sw(sw));
	wire signed[17:0] vwire_7_37;
	reg signed[17:0] vreg_7_37;
	node n7_37(.left(vreg_6_37), .right(vreg_8_37), .up(vreg_7_38), .down(vreg_7_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_37), .sw(sw));
	wire signed[17:0] vwire_7_38;
	reg signed[17:0] vreg_7_38;
	node n7_38(.left(vreg_6_38), .right(vreg_8_38), .up(vreg_7_39), .down(vreg_7_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_38), .sw(sw));
	wire signed[17:0] vwire_7_39;
	reg signed[17:0] vreg_7_39;
	node n7_39(.left(vreg_6_39), .right(vreg_8_39), .up(vreg_7_40), .down(vreg_7_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_39), .sw(sw));
	wire signed[17:0] vwire_7_40;
	reg signed[17:0] vreg_7_40;
	node n7_40(.left(vreg_6_40), .right(vreg_8_40), .up(vreg_7_41), .down(vreg_7_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_40), .sw(sw));
	wire signed[17:0] vwire_7_41;
	reg signed[17:0] vreg_7_41;
	node n7_41(.left(vreg_6_41), .right(vreg_8_41), .up(vreg_7_42), .down(vreg_7_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_41), .sw(sw));
	wire signed[17:0] vwire_7_42;
	reg signed[17:0] vreg_7_42;
	node n7_42(.left(vreg_6_42), .right(vreg_8_42), .up(vreg_7_43), .down(vreg_7_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_42), .sw(sw));
	wire signed[17:0] vwire_7_43;
	reg signed[17:0] vreg_7_43;
	node n7_43(.left(vreg_6_43), .right(vreg_8_43), .up(vreg_7_44), .down(vreg_7_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_43), .sw(sw));
	wire signed[17:0] vwire_7_44;
	reg signed[17:0] vreg_7_44;
	node n7_44(.left(vreg_6_44), .right(vreg_8_44), .up(vreg_7_45), .down(vreg_7_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_44), .sw(sw));
	wire signed[17:0] vwire_7_45;
	reg signed[17:0] vreg_7_45;
	node n7_45(.left(vreg_6_45), .right(vreg_8_45), .up(vreg_7_46), .down(vreg_7_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_45), .sw(sw));
	wire signed[17:0] vwire_7_46;
	reg signed[17:0] vreg_7_46;
	node n7_46(.left(vreg_6_46), .right(vreg_8_46), .up(vreg_7_47), .down(vreg_7_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_46), .sw(sw));
	wire signed[17:0] vwire_7_47;
	reg signed[17:0] vreg_7_47;
	node n7_47(.left(vreg_6_47), .right(vreg_8_47), .up(vreg_7_48), .down(vreg_7_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_47), .sw(sw));
	wire signed[17:0] vwire_7_48;
	reg signed[17:0] vreg_7_48;
	node n7_48(.left(vreg_6_48), .right(vreg_8_48), .up(vreg_7_49), .down(vreg_7_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_48), .sw(sw));
	wire signed[17:0] vwire_7_49;
	reg signed[17:0] vreg_7_49;
	node n7_49(.left(vreg_6_49), .right(vreg_8_49), .up(18'b0), .down(vreg_7_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_49), .sw(sw));
	wire signed[17:0] vwire_8_0;
	reg signed[17:0] vreg_8_0;
	node n8_0(.left(vreg_7_0), .right(vreg_9_0), .up(vreg_8_1), .down(vreg_8_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_0), .sw(sw));
	wire signed[17:0] vwire_8_1;
	reg signed[17:0] vreg_8_1;
	node n8_1(.left(vreg_7_1), .right(vreg_9_1), .up(vreg_8_2), .down(vreg_8_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_1), .sw(sw));
	wire signed[17:0] vwire_8_2;
	reg signed[17:0] vreg_8_2;
	node n8_2(.left(vreg_7_2), .right(vreg_9_2), .up(vreg_8_3), .down(vreg_8_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_2), .sw(sw));
	wire signed[17:0] vwire_8_3;
	reg signed[17:0] vreg_8_3;
	node n8_3(.left(vreg_7_3), .right(vreg_9_3), .up(vreg_8_4), .down(vreg_8_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_3), .sw(sw));
	wire signed[17:0] vwire_8_4;
	reg signed[17:0] vreg_8_4;
	node n8_4(.left(vreg_7_4), .right(vreg_9_4), .up(vreg_8_5), .down(vreg_8_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_4), .sw(sw));
	wire signed[17:0] vwire_8_5;
	reg signed[17:0] vreg_8_5;
	node n8_5(.left(vreg_7_5), .right(vreg_9_5), .up(vreg_8_6), .down(vreg_8_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_5), .sw(sw));
	wire signed[17:0] vwire_8_6;
	reg signed[17:0] vreg_8_6;
	node n8_6(.left(vreg_7_6), .right(vreg_9_6), .up(vreg_8_7), .down(vreg_8_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_6), .sw(sw));
	wire signed[17:0] vwire_8_7;
	reg signed[17:0] vreg_8_7;
	node n8_7(.left(vreg_7_7), .right(vreg_9_7), .up(vreg_8_8), .down(vreg_8_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_7), .sw(sw));
	wire signed[17:0] vwire_8_8;
	reg signed[17:0] vreg_8_8;
	node n8_8(.left(vreg_7_8), .right(vreg_9_8), .up(vreg_8_9), .down(vreg_8_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_8), .sw(sw));
	wire signed[17:0] vwire_8_9;
	reg signed[17:0] vreg_8_9;
	node n8_9(.left(vreg_7_9), .right(vreg_9_9), .up(vreg_8_10), .down(vreg_8_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_9), .sw(sw));
	wire signed[17:0] vwire_8_10;
	reg signed[17:0] vreg_8_10;
	node n8_10(.left(vreg_7_10), .right(vreg_9_10), .up(vreg_8_11), .down(vreg_8_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_10), .sw(sw));
	wire signed[17:0] vwire_8_11;
	reg signed[17:0] vreg_8_11;
	node n8_11(.left(vreg_7_11), .right(vreg_9_11), .up(vreg_8_12), .down(vreg_8_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_11), .sw(sw));
	wire signed[17:0] vwire_8_12;
	reg signed[17:0] vreg_8_12;
	node n8_12(.left(vreg_7_12), .right(vreg_9_12), .up(vreg_8_13), .down(vreg_8_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_12), .sw(sw));
	wire signed[17:0] vwire_8_13;
	reg signed[17:0] vreg_8_13;
	node n8_13(.left(vreg_7_13), .right(vreg_9_13), .up(vreg_8_14), .down(vreg_8_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_13), .sw(sw));
	wire signed[17:0] vwire_8_14;
	reg signed[17:0] vreg_8_14;
	node n8_14(.left(vreg_7_14), .right(vreg_9_14), .up(vreg_8_15), .down(vreg_8_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_14), .sw(sw));
	wire signed[17:0] vwire_8_15;
	reg signed[17:0] vreg_8_15;
	node n8_15(.left(vreg_7_15), .right(vreg_9_15), .up(vreg_8_16), .down(vreg_8_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_15), .sw(sw));
	wire signed[17:0] vwire_8_16;
	reg signed[17:0] vreg_8_16;
	node n8_16(.left(vreg_7_16), .right(vreg_9_16), .up(vreg_8_17), .down(vreg_8_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_16), .sw(sw));
	wire signed[17:0] vwire_8_17;
	reg signed[17:0] vreg_8_17;
	node n8_17(.left(vreg_7_17), .right(vreg_9_17), .up(vreg_8_18), .down(vreg_8_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_17), .sw(sw));
	wire signed[17:0] vwire_8_18;
	reg signed[17:0] vreg_8_18;
	node n8_18(.left(vreg_7_18), .right(vreg_9_18), .up(vreg_8_19), .down(vreg_8_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_18), .sw(sw));
	wire signed[17:0] vwire_8_19;
	reg signed[17:0] vreg_8_19;
	node n8_19(.left(vreg_7_19), .right(vreg_9_19), .up(vreg_8_20), .down(vreg_8_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_19), .sw(sw));
	wire signed[17:0] vwire_8_20;
	reg signed[17:0] vreg_8_20;
	node n8_20(.left(vreg_7_20), .right(vreg_9_20), .up(vreg_8_21), .down(vreg_8_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_20), .sw(sw));
	wire signed[17:0] vwire_8_21;
	reg signed[17:0] vreg_8_21;
	node n8_21(.left(vreg_7_21), .right(vreg_9_21), .up(vreg_8_22), .down(vreg_8_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_21), .sw(sw));
	wire signed[17:0] vwire_8_22;
	reg signed[17:0] vreg_8_22;
	node n8_22(.left(vreg_7_22), .right(vreg_9_22), .up(vreg_8_23), .down(vreg_8_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_22), .sw(sw));
	wire signed[17:0] vwire_8_23;
	reg signed[17:0] vreg_8_23;
	node n8_23(.left(vreg_7_23), .right(vreg_9_23), .up(vreg_8_24), .down(vreg_8_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_23), .sw(sw));
	wire signed[17:0] vwire_8_24;
	reg signed[17:0] vreg_8_24;
	node n8_24(.left(vreg_7_24), .right(vreg_9_24), .up(vreg_8_25), .down(vreg_8_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_24), .sw(sw));
	wire signed[17:0] vwire_8_25;
	reg signed[17:0] vreg_8_25;
	node n8_25(.left(vreg_7_25), .right(vreg_9_25), .up(vreg_8_26), .down(vreg_8_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_25), .sw(sw));
	wire signed[17:0] vwire_8_26;
	reg signed[17:0] vreg_8_26;
	node n8_26(.left(vreg_7_26), .right(vreg_9_26), .up(vreg_8_27), .down(vreg_8_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_26), .sw(sw));
	wire signed[17:0] vwire_8_27;
	reg signed[17:0] vreg_8_27;
	node n8_27(.left(vreg_7_27), .right(vreg_9_27), .up(vreg_8_28), .down(vreg_8_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_27), .sw(sw));
	wire signed[17:0] vwire_8_28;
	reg signed[17:0] vreg_8_28;
	node n8_28(.left(vreg_7_28), .right(vreg_9_28), .up(vreg_8_29), .down(vreg_8_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_28), .sw(sw));
	wire signed[17:0] vwire_8_29;
	reg signed[17:0] vreg_8_29;
	node n8_29(.left(vreg_7_29), .right(vreg_9_29), .up(vreg_8_30), .down(vreg_8_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_29), .sw(sw));
	wire signed[17:0] vwire_8_30;
	reg signed[17:0] vreg_8_30;
	node n8_30(.left(vreg_7_30), .right(vreg_9_30), .up(vreg_8_31), .down(vreg_8_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_30), .sw(sw));
	wire signed[17:0] vwire_8_31;
	reg signed[17:0] vreg_8_31;
	node n8_31(.left(vreg_7_31), .right(vreg_9_31), .up(vreg_8_32), .down(vreg_8_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_31), .sw(sw));
	wire signed[17:0] vwire_8_32;
	reg signed[17:0] vreg_8_32;
	node n8_32(.left(vreg_7_32), .right(vreg_9_32), .up(vreg_8_33), .down(vreg_8_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_32), .sw(sw));
	wire signed[17:0] vwire_8_33;
	reg signed[17:0] vreg_8_33;
	node n8_33(.left(vreg_7_33), .right(vreg_9_33), .up(vreg_8_34), .down(vreg_8_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_33), .sw(sw));
	wire signed[17:0] vwire_8_34;
	reg signed[17:0] vreg_8_34;
	node n8_34(.left(vreg_7_34), .right(vreg_9_34), .up(vreg_8_35), .down(vreg_8_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_34), .sw(sw));
	wire signed[17:0] vwire_8_35;
	reg signed[17:0] vreg_8_35;
	node n8_35(.left(vreg_7_35), .right(vreg_9_35), .up(vreg_8_36), .down(vreg_8_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_35), .sw(sw));
	wire signed[17:0] vwire_8_36;
	reg signed[17:0] vreg_8_36;
	node n8_36(.left(vreg_7_36), .right(vreg_9_36), .up(vreg_8_37), .down(vreg_8_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_36), .sw(sw));
	wire signed[17:0] vwire_8_37;
	reg signed[17:0] vreg_8_37;
	node n8_37(.left(vreg_7_37), .right(vreg_9_37), .up(vreg_8_38), .down(vreg_8_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_37), .sw(sw));
	wire signed[17:0] vwire_8_38;
	reg signed[17:0] vreg_8_38;
	node n8_38(.left(vreg_7_38), .right(vreg_9_38), .up(vreg_8_39), .down(vreg_8_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_38), .sw(sw));
	wire signed[17:0] vwire_8_39;
	reg signed[17:0] vreg_8_39;
	node n8_39(.left(vreg_7_39), .right(vreg_9_39), .up(vreg_8_40), .down(vreg_8_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_39), .sw(sw));
	wire signed[17:0] vwire_8_40;
	reg signed[17:0] vreg_8_40;
	node n8_40(.left(vreg_7_40), .right(vreg_9_40), .up(vreg_8_41), .down(vreg_8_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_40), .sw(sw));
	wire signed[17:0] vwire_8_41;
	reg signed[17:0] vreg_8_41;
	node n8_41(.left(vreg_7_41), .right(vreg_9_41), .up(vreg_8_42), .down(vreg_8_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_41), .sw(sw));
	wire signed[17:0] vwire_8_42;
	reg signed[17:0] vreg_8_42;
	node n8_42(.left(vreg_7_42), .right(vreg_9_42), .up(vreg_8_43), .down(vreg_8_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_42), .sw(sw));
	wire signed[17:0] vwire_8_43;
	reg signed[17:0] vreg_8_43;
	node n8_43(.left(vreg_7_43), .right(vreg_9_43), .up(vreg_8_44), .down(vreg_8_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_43), .sw(sw));
	wire signed[17:0] vwire_8_44;
	reg signed[17:0] vreg_8_44;
	node n8_44(.left(vreg_7_44), .right(vreg_9_44), .up(vreg_8_45), .down(vreg_8_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_44), .sw(sw));
	wire signed[17:0] vwire_8_45;
	reg signed[17:0] vreg_8_45;
	node n8_45(.left(vreg_7_45), .right(vreg_9_45), .up(vreg_8_46), .down(vreg_8_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_45), .sw(sw));
	wire signed[17:0] vwire_8_46;
	reg signed[17:0] vreg_8_46;
	node n8_46(.left(vreg_7_46), .right(vreg_9_46), .up(vreg_8_47), .down(vreg_8_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_46), .sw(sw));
	wire signed[17:0] vwire_8_47;
	reg signed[17:0] vreg_8_47;
	node n8_47(.left(vreg_7_47), .right(vreg_9_47), .up(vreg_8_48), .down(vreg_8_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_47), .sw(sw));
	wire signed[17:0] vwire_8_48;
	reg signed[17:0] vreg_8_48;
	node n8_48(.left(vreg_7_48), .right(vreg_9_48), .up(vreg_8_49), .down(vreg_8_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_48), .sw(sw));
	wire signed[17:0] vwire_8_49;
	reg signed[17:0] vreg_8_49;
	node n8_49(.left(vreg_7_49), .right(vreg_9_49), .up(18'b0), .down(vreg_8_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_8_49), .sw(sw));
	wire signed[17:0] vwire_9_0;
	reg signed[17:0] vreg_9_0;
	node n9_0(.left(vreg_8_0), .right(vreg_10_0), .up(vreg_9_1), .down(vreg_9_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_0), .sw(sw));
	wire signed[17:0] vwire_9_1;
	reg signed[17:0] vreg_9_1;
	node n9_1(.left(vreg_8_1), .right(vreg_10_1), .up(vreg_9_2), .down(vreg_9_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_1), .sw(sw));
	wire signed[17:0] vwire_9_2;
	reg signed[17:0] vreg_9_2;
	node n9_2(.left(vreg_8_2), .right(vreg_10_2), .up(vreg_9_3), .down(vreg_9_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_2), .sw(sw));
	wire signed[17:0] vwire_9_3;
	reg signed[17:0] vreg_9_3;
	node n9_3(.left(vreg_8_3), .right(vreg_10_3), .up(vreg_9_4), .down(vreg_9_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_3), .sw(sw));
	wire signed[17:0] vwire_9_4;
	reg signed[17:0] vreg_9_4;
	node n9_4(.left(vreg_8_4), .right(vreg_10_4), .up(vreg_9_5), .down(vreg_9_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_4), .sw(sw));
	wire signed[17:0] vwire_9_5;
	reg signed[17:0] vreg_9_5;
	node n9_5(.left(vreg_8_5), .right(vreg_10_5), .up(vreg_9_6), .down(vreg_9_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_5), .sw(sw));
	wire signed[17:0] vwire_9_6;
	reg signed[17:0] vreg_9_6;
	node n9_6(.left(vreg_8_6), .right(vreg_10_6), .up(vreg_9_7), .down(vreg_9_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_6), .sw(sw));
	wire signed[17:0] vwire_9_7;
	reg signed[17:0] vreg_9_7;
	node n9_7(.left(vreg_8_7), .right(vreg_10_7), .up(vreg_9_8), .down(vreg_9_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_7), .sw(sw));
	wire signed[17:0] vwire_9_8;
	reg signed[17:0] vreg_9_8;
	node n9_8(.left(vreg_8_8), .right(vreg_10_8), .up(vreg_9_9), .down(vreg_9_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_8), .sw(sw));
	wire signed[17:0] vwire_9_9;
	reg signed[17:0] vreg_9_9;
	node n9_9(.left(vreg_8_9), .right(vreg_10_9), .up(vreg_9_10), .down(vreg_9_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_9), .sw(sw));
	wire signed[17:0] vwire_9_10;
	reg signed[17:0] vreg_9_10;
	node n9_10(.left(vreg_8_10), .right(vreg_10_10), .up(vreg_9_11), .down(vreg_9_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_10), .sw(sw));
	wire signed[17:0] vwire_9_11;
	reg signed[17:0] vreg_9_11;
	node n9_11(.left(vreg_8_11), .right(vreg_10_11), .up(vreg_9_12), .down(vreg_9_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_11), .sw(sw));
	wire signed[17:0] vwire_9_12;
	reg signed[17:0] vreg_9_12;
	node n9_12(.left(vreg_8_12), .right(vreg_10_12), .up(vreg_9_13), .down(vreg_9_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_12), .sw(sw));
	wire signed[17:0] vwire_9_13;
	reg signed[17:0] vreg_9_13;
	node n9_13(.left(vreg_8_13), .right(vreg_10_13), .up(vreg_9_14), .down(vreg_9_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_13), .sw(sw));
	wire signed[17:0] vwire_9_14;
	reg signed[17:0] vreg_9_14;
	node n9_14(.left(vreg_8_14), .right(vreg_10_14), .up(vreg_9_15), .down(vreg_9_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_14), .sw(sw));
	wire signed[17:0] vwire_9_15;
	reg signed[17:0] vreg_9_15;
	node n9_15(.left(vreg_8_15), .right(vreg_10_15), .up(vreg_9_16), .down(vreg_9_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_15), .sw(sw));
	wire signed[17:0] vwire_9_16;
	reg signed[17:0] vreg_9_16;
	node n9_16(.left(vreg_8_16), .right(vreg_10_16), .up(vreg_9_17), .down(vreg_9_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_16), .sw(sw));
	wire signed[17:0] vwire_9_17;
	reg signed[17:0] vreg_9_17;
	node n9_17(.left(vreg_8_17), .right(vreg_10_17), .up(vreg_9_18), .down(vreg_9_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_17), .sw(sw));
	wire signed[17:0] vwire_9_18;
	reg signed[17:0] vreg_9_18;
	node n9_18(.left(vreg_8_18), .right(vreg_10_18), .up(vreg_9_19), .down(vreg_9_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_18), .sw(sw));
	wire signed[17:0] vwire_9_19;
	reg signed[17:0] vreg_9_19;
	node n9_19(.left(vreg_8_19), .right(vreg_10_19), .up(vreg_9_20), .down(vreg_9_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_19), .sw(sw));
	wire signed[17:0] vwire_9_20;
	reg signed[17:0] vreg_9_20;
	node n9_20(.left(vreg_8_20), .right(vreg_10_20), .up(vreg_9_21), .down(vreg_9_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_20), .sw(sw));
	wire signed[17:0] vwire_9_21;
	reg signed[17:0] vreg_9_21;
	node n9_21(.left(vreg_8_21), .right(vreg_10_21), .up(vreg_9_22), .down(vreg_9_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_21), .sw(sw));
	wire signed[17:0] vwire_9_22;
	reg signed[17:0] vreg_9_22;
	node n9_22(.left(vreg_8_22), .right(vreg_10_22), .up(vreg_9_23), .down(vreg_9_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_22), .sw(sw));
	wire signed[17:0] vwire_9_23;
	reg signed[17:0] vreg_9_23;
	node n9_23(.left(vreg_8_23), .right(vreg_10_23), .up(vreg_9_24), .down(vreg_9_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_23), .sw(sw));
	wire signed[17:0] vwire_9_24;
	reg signed[17:0] vreg_9_24;
	node n9_24(.left(vreg_8_24), .right(vreg_10_24), .up(vreg_9_25), .down(vreg_9_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_24), .sw(sw));
	wire signed[17:0] vwire_9_25;
	reg signed[17:0] vreg_9_25;
	node n9_25(.left(vreg_8_25), .right(vreg_10_25), .up(vreg_9_26), .down(vreg_9_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_25), .sw(sw));
	wire signed[17:0] vwire_9_26;
	reg signed[17:0] vreg_9_26;
	node n9_26(.left(vreg_8_26), .right(vreg_10_26), .up(vreg_9_27), .down(vreg_9_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_26), .sw(sw));
	wire signed[17:0] vwire_9_27;
	reg signed[17:0] vreg_9_27;
	node n9_27(.left(vreg_8_27), .right(vreg_10_27), .up(vreg_9_28), .down(vreg_9_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_27), .sw(sw));
	wire signed[17:0] vwire_9_28;
	reg signed[17:0] vreg_9_28;
	node n9_28(.left(vreg_8_28), .right(vreg_10_28), .up(vreg_9_29), .down(vreg_9_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_28), .sw(sw));
	wire signed[17:0] vwire_9_29;
	reg signed[17:0] vreg_9_29;
	node n9_29(.left(vreg_8_29), .right(vreg_10_29), .up(vreg_9_30), .down(vreg_9_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_29), .sw(sw));
	wire signed[17:0] vwire_9_30;
	reg signed[17:0] vreg_9_30;
	node n9_30(.left(vreg_8_30), .right(vreg_10_30), .up(vreg_9_31), .down(vreg_9_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_30), .sw(sw));
	wire signed[17:0] vwire_9_31;
	reg signed[17:0] vreg_9_31;
	node n9_31(.left(vreg_8_31), .right(vreg_10_31), .up(vreg_9_32), .down(vreg_9_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_31), .sw(sw));
	wire signed[17:0] vwire_9_32;
	reg signed[17:0] vreg_9_32;
	node n9_32(.left(vreg_8_32), .right(vreg_10_32), .up(vreg_9_33), .down(vreg_9_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_32), .sw(sw));
	wire signed[17:0] vwire_9_33;
	reg signed[17:0] vreg_9_33;
	node n9_33(.left(vreg_8_33), .right(vreg_10_33), .up(vreg_9_34), .down(vreg_9_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_33), .sw(sw));
	wire signed[17:0] vwire_9_34;
	reg signed[17:0] vreg_9_34;
	node n9_34(.left(vreg_8_34), .right(vreg_10_34), .up(vreg_9_35), .down(vreg_9_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_34), .sw(sw));
	wire signed[17:0] vwire_9_35;
	reg signed[17:0] vreg_9_35;
	node n9_35(.left(vreg_8_35), .right(vreg_10_35), .up(vreg_9_36), .down(vreg_9_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_35), .sw(sw));
	wire signed[17:0] vwire_9_36;
	reg signed[17:0] vreg_9_36;
	node n9_36(.left(vreg_8_36), .right(vreg_10_36), .up(vreg_9_37), .down(vreg_9_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_36), .sw(sw));
	wire signed[17:0] vwire_9_37;
	reg signed[17:0] vreg_9_37;
	node n9_37(.left(vreg_8_37), .right(vreg_10_37), .up(vreg_9_38), .down(vreg_9_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_37), .sw(sw));
	wire signed[17:0] vwire_9_38;
	reg signed[17:0] vreg_9_38;
	node n9_38(.left(vreg_8_38), .right(vreg_10_38), .up(vreg_9_39), .down(vreg_9_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_38), .sw(sw));
	wire signed[17:0] vwire_9_39;
	reg signed[17:0] vreg_9_39;
	node n9_39(.left(vreg_8_39), .right(vreg_10_39), .up(vreg_9_40), .down(vreg_9_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_39), .sw(sw));
	wire signed[17:0] vwire_9_40;
	reg signed[17:0] vreg_9_40;
	node n9_40(.left(vreg_8_40), .right(vreg_10_40), .up(vreg_9_41), .down(vreg_9_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_40), .sw(sw));
	wire signed[17:0] vwire_9_41;
	reg signed[17:0] vreg_9_41;
	node n9_41(.left(vreg_8_41), .right(vreg_10_41), .up(vreg_9_42), .down(vreg_9_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_41), .sw(sw));
	wire signed[17:0] vwire_9_42;
	reg signed[17:0] vreg_9_42;
	node n9_42(.left(vreg_8_42), .right(vreg_10_42), .up(vreg_9_43), .down(vreg_9_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_42), .sw(sw));
	wire signed[17:0] vwire_9_43;
	reg signed[17:0] vreg_9_43;
	node n9_43(.left(vreg_8_43), .right(vreg_10_43), .up(vreg_9_44), .down(vreg_9_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_43), .sw(sw));
	wire signed[17:0] vwire_9_44;
	reg signed[17:0] vreg_9_44;
	node n9_44(.left(vreg_8_44), .right(vreg_10_44), .up(vreg_9_45), .down(vreg_9_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_44), .sw(sw));
	wire signed[17:0] vwire_9_45;
	reg signed[17:0] vreg_9_45;
	node n9_45(.left(vreg_8_45), .right(vreg_10_45), .up(vreg_9_46), .down(vreg_9_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_45), .sw(sw));
	wire signed[17:0] vwire_9_46;
	reg signed[17:0] vreg_9_46;
	node n9_46(.left(vreg_8_46), .right(vreg_10_46), .up(vreg_9_47), .down(vreg_9_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_46), .sw(sw));
	wire signed[17:0] vwire_9_47;
	reg signed[17:0] vreg_9_47;
	node n9_47(.left(vreg_8_47), .right(vreg_10_47), .up(vreg_9_48), .down(vreg_9_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_47), .sw(sw));
	wire signed[17:0] vwire_9_48;
	reg signed[17:0] vreg_9_48;
	node n9_48(.left(vreg_8_48), .right(vreg_10_48), .up(vreg_9_49), .down(vreg_9_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_48), .sw(sw));
	wire signed[17:0] vwire_9_49;
	reg signed[17:0] vreg_9_49;
	node n9_49(.left(vreg_8_49), .right(vreg_10_49), .up(18'b0), .down(vreg_9_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_9_49), .sw(sw));
	wire signed[17:0] vwire_10_0;
	reg signed[17:0] vreg_10_0;
	node n10_0(.left(vreg_9_0), .right(vreg_11_0), .up(vreg_10_1), .down(vreg_10_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_0), .sw(sw));
	wire signed[17:0] vwire_10_1;
	reg signed[17:0] vreg_10_1;
	node n10_1(.left(vreg_9_1), .right(vreg_11_1), .up(vreg_10_2), .down(vreg_10_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_1), .sw(sw));
	wire signed[17:0] vwire_10_2;
	reg signed[17:0] vreg_10_2;
	node n10_2(.left(vreg_9_2), .right(vreg_11_2), .up(vreg_10_3), .down(vreg_10_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_2), .sw(sw));
	wire signed[17:0] vwire_10_3;
	reg signed[17:0] vreg_10_3;
	node n10_3(.left(vreg_9_3), .right(vreg_11_3), .up(vreg_10_4), .down(vreg_10_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_3), .sw(sw));
	wire signed[17:0] vwire_10_4;
	reg signed[17:0] vreg_10_4;
	node n10_4(.left(vreg_9_4), .right(vreg_11_4), .up(vreg_10_5), .down(vreg_10_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_4), .sw(sw));
	wire signed[17:0] vwire_10_5;
	reg signed[17:0] vreg_10_5;
	node n10_5(.left(vreg_9_5), .right(vreg_11_5), .up(vreg_10_6), .down(vreg_10_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_5), .sw(sw));
	wire signed[17:0] vwire_10_6;
	reg signed[17:0] vreg_10_6;
	node n10_6(.left(vreg_9_6), .right(vreg_11_6), .up(vreg_10_7), .down(vreg_10_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_6), .sw(sw));
	wire signed[17:0] vwire_10_7;
	reg signed[17:0] vreg_10_7;
	node n10_7(.left(vreg_9_7), .right(vreg_11_7), .up(vreg_10_8), .down(vreg_10_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_7), .sw(sw));
	wire signed[17:0] vwire_10_8;
	reg signed[17:0] vreg_10_8;
	node n10_8(.left(vreg_9_8), .right(vreg_11_8), .up(vreg_10_9), .down(vreg_10_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_8), .sw(sw));
	wire signed[17:0] vwire_10_9;
	reg signed[17:0] vreg_10_9;
	node n10_9(.left(vreg_9_9), .right(vreg_11_9), .up(vreg_10_10), .down(vreg_10_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_9), .sw(sw));
	wire signed[17:0] vwire_10_10;
	reg signed[17:0] vreg_10_10;
	node n10_10(.left(vreg_9_10), .right(vreg_11_10), .up(vreg_10_11), .down(vreg_10_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_10), .sw(sw));
	wire signed[17:0] vwire_10_11;
	reg signed[17:0] vreg_10_11;
	node n10_11(.left(vreg_9_11), .right(vreg_11_11), .up(vreg_10_12), .down(vreg_10_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_11), .sw(sw));
	wire signed[17:0] vwire_10_12;
	reg signed[17:0] vreg_10_12;
	node n10_12(.left(vreg_9_12), .right(vreg_11_12), .up(vreg_10_13), .down(vreg_10_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_12), .sw(sw));
	wire signed[17:0] vwire_10_13;
	reg signed[17:0] vreg_10_13;
	node n10_13(.left(vreg_9_13), .right(vreg_11_13), .up(vreg_10_14), .down(vreg_10_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_13), .sw(sw));
	wire signed[17:0] vwire_10_14;
	reg signed[17:0] vreg_10_14;
	node n10_14(.left(vreg_9_14), .right(vreg_11_14), .up(vreg_10_15), .down(vreg_10_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_14), .sw(sw));
	wire signed[17:0] vwire_10_15;
	reg signed[17:0] vreg_10_15;
	node n10_15(.left(vreg_9_15), .right(vreg_11_15), .up(vreg_10_16), .down(vreg_10_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_15), .sw(sw));
	wire signed[17:0] vwire_10_16;
	reg signed[17:0] vreg_10_16;
	node n10_16(.left(vreg_9_16), .right(vreg_11_16), .up(vreg_10_17), .down(vreg_10_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_16), .sw(sw));
	wire signed[17:0] vwire_10_17;
	reg signed[17:0] vreg_10_17;
	node n10_17(.left(vreg_9_17), .right(vreg_11_17), .up(vreg_10_18), .down(vreg_10_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_17), .sw(sw));
	wire signed[17:0] vwire_10_18;
	reg signed[17:0] vreg_10_18;
	node n10_18(.left(vreg_9_18), .right(vreg_11_18), .up(vreg_10_19), .down(vreg_10_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_18), .sw(sw));
	wire signed[17:0] vwire_10_19;
	reg signed[17:0] vreg_10_19;
	node n10_19(.left(vreg_9_19), .right(vreg_11_19), .up(vreg_10_20), .down(vreg_10_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_19), .sw(sw));
	wire signed[17:0] vwire_10_20;
	reg signed[17:0] vreg_10_20;
	node n10_20(.left(vreg_9_20), .right(vreg_11_20), .up(vreg_10_21), .down(vreg_10_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_20), .sw(sw));
	wire signed[17:0] vwire_10_21;
	reg signed[17:0] vreg_10_21;
	node n10_21(.left(vreg_9_21), .right(vreg_11_21), .up(vreg_10_22), .down(vreg_10_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_21), .sw(sw));
	wire signed[17:0] vwire_10_22;
	reg signed[17:0] vreg_10_22;
	node n10_22(.left(vreg_9_22), .right(vreg_11_22), .up(vreg_10_23), .down(vreg_10_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_22), .sw(sw));
	wire signed[17:0] vwire_10_23;
	reg signed[17:0] vreg_10_23;
	node n10_23(.left(vreg_9_23), .right(vreg_11_23), .up(vreg_10_24), .down(vreg_10_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_23), .sw(sw));
	wire signed[17:0] vwire_10_24;
	reg signed[17:0] vreg_10_24;
	node n10_24(.left(vreg_9_24), .right(vreg_11_24), .up(vreg_10_25), .down(vreg_10_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_24), .sw(sw));
	wire signed[17:0] vwire_10_25;
	reg signed[17:0] vreg_10_25;
	node n10_25(.left(vreg_9_25), .right(vreg_11_25), .up(vreg_10_26), .down(vreg_10_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_25), .sw(sw));
	wire signed[17:0] vwire_10_26;
	reg signed[17:0] vreg_10_26;
	node n10_26(.left(vreg_9_26), .right(vreg_11_26), .up(vreg_10_27), .down(vreg_10_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_26), .sw(sw));
	wire signed[17:0] vwire_10_27;
	reg signed[17:0] vreg_10_27;
	node n10_27(.left(vreg_9_27), .right(vreg_11_27), .up(vreg_10_28), .down(vreg_10_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_27), .sw(sw));
	wire signed[17:0] vwire_10_28;
	reg signed[17:0] vreg_10_28;
	node n10_28(.left(vreg_9_28), .right(vreg_11_28), .up(vreg_10_29), .down(vreg_10_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_28), .sw(sw));
	wire signed[17:0] vwire_10_29;
	reg signed[17:0] vreg_10_29;
	node n10_29(.left(vreg_9_29), .right(vreg_11_29), .up(vreg_10_30), .down(vreg_10_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_29), .sw(sw));
	wire signed[17:0] vwire_10_30;
	reg signed[17:0] vreg_10_30;
	node n10_30(.left(vreg_9_30), .right(vreg_11_30), .up(vreg_10_31), .down(vreg_10_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_30), .sw(sw));
	wire signed[17:0] vwire_10_31;
	reg signed[17:0] vreg_10_31;
	node n10_31(.left(vreg_9_31), .right(vreg_11_31), .up(vreg_10_32), .down(vreg_10_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_31), .sw(sw));
	wire signed[17:0] vwire_10_32;
	reg signed[17:0] vreg_10_32;
	node n10_32(.left(vreg_9_32), .right(vreg_11_32), .up(vreg_10_33), .down(vreg_10_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_32), .sw(sw));
	wire signed[17:0] vwire_10_33;
	reg signed[17:0] vreg_10_33;
	node n10_33(.left(vreg_9_33), .right(vreg_11_33), .up(vreg_10_34), .down(vreg_10_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_33), .sw(sw));
	wire signed[17:0] vwire_10_34;
	reg signed[17:0] vreg_10_34;
	node n10_34(.left(vreg_9_34), .right(vreg_11_34), .up(vreg_10_35), .down(vreg_10_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_34), .sw(sw));
	wire signed[17:0] vwire_10_35;
	reg signed[17:0] vreg_10_35;
	node n10_35(.left(vreg_9_35), .right(vreg_11_35), .up(vreg_10_36), .down(vreg_10_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_35), .sw(sw));
	wire signed[17:0] vwire_10_36;
	reg signed[17:0] vreg_10_36;
	node n10_36(.left(vreg_9_36), .right(vreg_11_36), .up(vreg_10_37), .down(vreg_10_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_36), .sw(sw));
	wire signed[17:0] vwire_10_37;
	reg signed[17:0] vreg_10_37;
	node n10_37(.left(vreg_9_37), .right(vreg_11_37), .up(vreg_10_38), .down(vreg_10_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_37), .sw(sw));
	wire signed[17:0] vwire_10_38;
	reg signed[17:0] vreg_10_38;
	node n10_38(.left(vreg_9_38), .right(vreg_11_38), .up(vreg_10_39), .down(vreg_10_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_38), .sw(sw));
	wire signed[17:0] vwire_10_39;
	reg signed[17:0] vreg_10_39;
	node n10_39(.left(vreg_9_39), .right(vreg_11_39), .up(vreg_10_40), .down(vreg_10_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_39), .sw(sw));
	wire signed[17:0] vwire_10_40;
	reg signed[17:0] vreg_10_40;
	node n10_40(.left(vreg_9_40), .right(vreg_11_40), .up(vreg_10_41), .down(vreg_10_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_40), .sw(sw));
	wire signed[17:0] vwire_10_41;
	reg signed[17:0] vreg_10_41;
	node n10_41(.left(vreg_9_41), .right(vreg_11_41), .up(vreg_10_42), .down(vreg_10_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_41), .sw(sw));
	wire signed[17:0] vwire_10_42;
	reg signed[17:0] vreg_10_42;
	node n10_42(.left(vreg_9_42), .right(vreg_11_42), .up(vreg_10_43), .down(vreg_10_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_42), .sw(sw));
	wire signed[17:0] vwire_10_43;
	reg signed[17:0] vreg_10_43;
	node n10_43(.left(vreg_9_43), .right(vreg_11_43), .up(vreg_10_44), .down(vreg_10_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_43), .sw(sw));
	wire signed[17:0] vwire_10_44;
	reg signed[17:0] vreg_10_44;
	node n10_44(.left(vreg_9_44), .right(vreg_11_44), .up(vreg_10_45), .down(vreg_10_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_44), .sw(sw));
	wire signed[17:0] vwire_10_45;
	reg signed[17:0] vreg_10_45;
	node n10_45(.left(vreg_9_45), .right(vreg_11_45), .up(vreg_10_46), .down(vreg_10_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_45), .sw(sw));
	wire signed[17:0] vwire_10_46;
	reg signed[17:0] vreg_10_46;
	node n10_46(.left(vreg_9_46), .right(vreg_11_46), .up(vreg_10_47), .down(vreg_10_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_46), .sw(sw));
	wire signed[17:0] vwire_10_47;
	reg signed[17:0] vreg_10_47;
	node n10_47(.left(vreg_9_47), .right(vreg_11_47), .up(vreg_10_48), .down(vreg_10_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_47), .sw(sw));
	wire signed[17:0] vwire_10_48;
	reg signed[17:0] vreg_10_48;
	node n10_48(.left(vreg_9_48), .right(vreg_11_48), .up(vreg_10_49), .down(vreg_10_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_48), .sw(sw));
	wire signed[17:0] vwire_10_49;
	reg signed[17:0] vreg_10_49;
	node n10_49(.left(vreg_9_49), .right(vreg_11_49), .up(18'b0), .down(vreg_10_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_10_49), .sw(sw));
	wire signed[17:0] vwire_11_0;
	reg signed[17:0] vreg_11_0;
	node n11_0(.left(vreg_10_0), .right(vreg_12_0), .up(vreg_11_1), .down(vreg_11_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_0), .sw(sw));
	wire signed[17:0] vwire_11_1;
	reg signed[17:0] vreg_11_1;
	node n11_1(.left(vreg_10_1), .right(vreg_12_1), .up(vreg_11_2), .down(vreg_11_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_1), .sw(sw));
	wire signed[17:0] vwire_11_2;
	reg signed[17:0] vreg_11_2;
	node n11_2(.left(vreg_10_2), .right(vreg_12_2), .up(vreg_11_3), .down(vreg_11_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_2), .sw(sw));
	wire signed[17:0] vwire_11_3;
	reg signed[17:0] vreg_11_3;
	node n11_3(.left(vreg_10_3), .right(vreg_12_3), .up(vreg_11_4), .down(vreg_11_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_3), .sw(sw));
	wire signed[17:0] vwire_11_4;
	reg signed[17:0] vreg_11_4;
	node n11_4(.left(vreg_10_4), .right(vreg_12_4), .up(vreg_11_5), .down(vreg_11_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_4), .sw(sw));
	wire signed[17:0] vwire_11_5;
	reg signed[17:0] vreg_11_5;
	node n11_5(.left(vreg_10_5), .right(vreg_12_5), .up(vreg_11_6), .down(vreg_11_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_5), .sw(sw));
	wire signed[17:0] vwire_11_6;
	reg signed[17:0] vreg_11_6;
	node n11_6(.left(vreg_10_6), .right(vreg_12_6), .up(vreg_11_7), .down(vreg_11_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_6), .sw(sw));
	wire signed[17:0] vwire_11_7;
	reg signed[17:0] vreg_11_7;
	node n11_7(.left(vreg_10_7), .right(vreg_12_7), .up(vreg_11_8), .down(vreg_11_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_7), .sw(sw));
	wire signed[17:0] vwire_11_8;
	reg signed[17:0] vreg_11_8;
	node n11_8(.left(vreg_10_8), .right(vreg_12_8), .up(vreg_11_9), .down(vreg_11_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_8), .sw(sw));
	wire signed[17:0] vwire_11_9;
	reg signed[17:0] vreg_11_9;
	node n11_9(.left(vreg_10_9), .right(vreg_12_9), .up(vreg_11_10), .down(vreg_11_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_9), .sw(sw));
	wire signed[17:0] vwire_11_10;
	reg signed[17:0] vreg_11_10;
	node n11_10(.left(vreg_10_10), .right(vreg_12_10), .up(vreg_11_11), .down(vreg_11_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_10), .sw(sw));
	wire signed[17:0] vwire_11_11;
	reg signed[17:0] vreg_11_11;
	node n11_11(.left(vreg_10_11), .right(vreg_12_11), .up(vreg_11_12), .down(vreg_11_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_11), .sw(sw));
	wire signed[17:0] vwire_11_12;
	reg signed[17:0] vreg_11_12;
	node n11_12(.left(vreg_10_12), .right(vreg_12_12), .up(vreg_11_13), .down(vreg_11_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_12), .sw(sw));
	wire signed[17:0] vwire_11_13;
	reg signed[17:0] vreg_11_13;
	node n11_13(.left(vreg_10_13), .right(vreg_12_13), .up(vreg_11_14), .down(vreg_11_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_13), .sw(sw));
	wire signed[17:0] vwire_11_14;
	reg signed[17:0] vreg_11_14;
	node n11_14(.left(vreg_10_14), .right(vreg_12_14), .up(vreg_11_15), .down(vreg_11_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_14), .sw(sw));
	wire signed[17:0] vwire_11_15;
	reg signed[17:0] vreg_11_15;
	node n11_15(.left(vreg_10_15), .right(vreg_12_15), .up(vreg_11_16), .down(vreg_11_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_15), .sw(sw));
	wire signed[17:0] vwire_11_16;
	reg signed[17:0] vreg_11_16;
	node n11_16(.left(vreg_10_16), .right(vreg_12_16), .up(vreg_11_17), .down(vreg_11_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_16), .sw(sw));
	wire signed[17:0] vwire_11_17;
	reg signed[17:0] vreg_11_17;
	node n11_17(.left(vreg_10_17), .right(vreg_12_17), .up(vreg_11_18), .down(vreg_11_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_17), .sw(sw));
	wire signed[17:0] vwire_11_18;
	reg signed[17:0] vreg_11_18;
	node n11_18(.left(vreg_10_18), .right(vreg_12_18), .up(vreg_11_19), .down(vreg_11_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_18), .sw(sw));
	wire signed[17:0] vwire_11_19;
	reg signed[17:0] vreg_11_19;
	node n11_19(.left(vreg_10_19), .right(vreg_12_19), .up(vreg_11_20), .down(vreg_11_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_19), .sw(sw));
	wire signed[17:0] vwire_11_20;
	reg signed[17:0] vreg_11_20;
	node n11_20(.left(vreg_10_20), .right(vreg_12_20), .up(vreg_11_21), .down(vreg_11_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_20), .sw(sw));
	wire signed[17:0] vwire_11_21;
	reg signed[17:0] vreg_11_21;
	node n11_21(.left(vreg_10_21), .right(vreg_12_21), .up(vreg_11_22), .down(vreg_11_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_21), .sw(sw));
	wire signed[17:0] vwire_11_22;
	reg signed[17:0] vreg_11_22;
	node n11_22(.left(vreg_10_22), .right(vreg_12_22), .up(vreg_11_23), .down(vreg_11_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_22), .sw(sw));
	wire signed[17:0] vwire_11_23;
	reg signed[17:0] vreg_11_23;
	node n11_23(.left(vreg_10_23), .right(vreg_12_23), .up(vreg_11_24), .down(vreg_11_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_23), .sw(sw));
	wire signed[17:0] vwire_11_24;
	reg signed[17:0] vreg_11_24;
	node n11_24(.left(vreg_10_24), .right(vreg_12_24), .up(vreg_11_25), .down(vreg_11_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_24), .sw(sw));
	wire signed[17:0] vwire_11_25;
	reg signed[17:0] vreg_11_25;
	node n11_25(.left(vreg_10_25), .right(vreg_12_25), .up(vreg_11_26), .down(vreg_11_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_25), .sw(sw));
	wire signed[17:0] vwire_11_26;
	reg signed[17:0] vreg_11_26;
	node n11_26(.left(vreg_10_26), .right(vreg_12_26), .up(vreg_11_27), .down(vreg_11_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_26), .sw(sw));
	wire signed[17:0] vwire_11_27;
	reg signed[17:0] vreg_11_27;
	node n11_27(.left(vreg_10_27), .right(vreg_12_27), .up(vreg_11_28), .down(vreg_11_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_27), .sw(sw));
	wire signed[17:0] vwire_11_28;
	reg signed[17:0] vreg_11_28;
	node n11_28(.left(vreg_10_28), .right(vreg_12_28), .up(vreg_11_29), .down(vreg_11_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_28), .sw(sw));
	wire signed[17:0] vwire_11_29;
	reg signed[17:0] vreg_11_29;
	node n11_29(.left(vreg_10_29), .right(vreg_12_29), .up(vreg_11_30), .down(vreg_11_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_29), .sw(sw));
	wire signed[17:0] vwire_11_30;
	reg signed[17:0] vreg_11_30;
	node n11_30(.left(vreg_10_30), .right(vreg_12_30), .up(vreg_11_31), .down(vreg_11_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_30), .sw(sw));
	wire signed[17:0] vwire_11_31;
	reg signed[17:0] vreg_11_31;
	node n11_31(.left(vreg_10_31), .right(vreg_12_31), .up(vreg_11_32), .down(vreg_11_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_31), .sw(sw));
	wire signed[17:0] vwire_11_32;
	reg signed[17:0] vreg_11_32;
	node n11_32(.left(vreg_10_32), .right(vreg_12_32), .up(vreg_11_33), .down(vreg_11_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_32), .sw(sw));
	wire signed[17:0] vwire_11_33;
	reg signed[17:0] vreg_11_33;
	node n11_33(.left(vreg_10_33), .right(vreg_12_33), .up(vreg_11_34), .down(vreg_11_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_33), .sw(sw));
	wire signed[17:0] vwire_11_34;
	reg signed[17:0] vreg_11_34;
	node n11_34(.left(vreg_10_34), .right(vreg_12_34), .up(vreg_11_35), .down(vreg_11_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_34), .sw(sw));
	wire signed[17:0] vwire_11_35;
	reg signed[17:0] vreg_11_35;
	node n11_35(.left(vreg_10_35), .right(vreg_12_35), .up(vreg_11_36), .down(vreg_11_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_35), .sw(sw));
	wire signed[17:0] vwire_11_36;
	reg signed[17:0] vreg_11_36;
	node n11_36(.left(vreg_10_36), .right(vreg_12_36), .up(vreg_11_37), .down(vreg_11_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_36), .sw(sw));
	wire signed[17:0] vwire_11_37;
	reg signed[17:0] vreg_11_37;
	node n11_37(.left(vreg_10_37), .right(vreg_12_37), .up(vreg_11_38), .down(vreg_11_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_37), .sw(sw));
	wire signed[17:0] vwire_11_38;
	reg signed[17:0] vreg_11_38;
	node n11_38(.left(vreg_10_38), .right(vreg_12_38), .up(vreg_11_39), .down(vreg_11_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_38), .sw(sw));
	wire signed[17:0] vwire_11_39;
	reg signed[17:0] vreg_11_39;
	node n11_39(.left(vreg_10_39), .right(vreg_12_39), .up(vreg_11_40), .down(vreg_11_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_39), .sw(sw));
	wire signed[17:0] vwire_11_40;
	reg signed[17:0] vreg_11_40;
	node n11_40(.left(vreg_10_40), .right(vreg_12_40), .up(vreg_11_41), .down(vreg_11_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_40), .sw(sw));
	wire signed[17:0] vwire_11_41;
	reg signed[17:0] vreg_11_41;
	node n11_41(.left(vreg_10_41), .right(vreg_12_41), .up(vreg_11_42), .down(vreg_11_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_41), .sw(sw));
	wire signed[17:0] vwire_11_42;
	reg signed[17:0] vreg_11_42;
	node n11_42(.left(vreg_10_42), .right(vreg_12_42), .up(vreg_11_43), .down(vreg_11_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_42), .sw(sw));
	wire signed[17:0] vwire_11_43;
	reg signed[17:0] vreg_11_43;
	node n11_43(.left(vreg_10_43), .right(vreg_12_43), .up(vreg_11_44), .down(vreg_11_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_43), .sw(sw));
	wire signed[17:0] vwire_11_44;
	reg signed[17:0] vreg_11_44;
	node n11_44(.left(vreg_10_44), .right(vreg_12_44), .up(vreg_11_45), .down(vreg_11_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_44), .sw(sw));
	wire signed[17:0] vwire_11_45;
	reg signed[17:0] vreg_11_45;
	node n11_45(.left(vreg_10_45), .right(vreg_12_45), .up(vreg_11_46), .down(vreg_11_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_45), .sw(sw));
	wire signed[17:0] vwire_11_46;
	reg signed[17:0] vreg_11_46;
	node n11_46(.left(vreg_10_46), .right(vreg_12_46), .up(vreg_11_47), .down(vreg_11_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_46), .sw(sw));
	wire signed[17:0] vwire_11_47;
	reg signed[17:0] vreg_11_47;
	node n11_47(.left(vreg_10_47), .right(vreg_12_47), .up(vreg_11_48), .down(vreg_11_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_47), .sw(sw));
	wire signed[17:0] vwire_11_48;
	reg signed[17:0] vreg_11_48;
	node n11_48(.left(vreg_10_48), .right(vreg_12_48), .up(vreg_11_49), .down(vreg_11_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_48), .sw(sw));
	wire signed[17:0] vwire_11_49;
	reg signed[17:0] vreg_11_49;
	node n11_49(.left(vreg_10_49), .right(vreg_12_49), .up(18'b0), .down(vreg_11_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_11_49), .sw(sw));
	wire signed[17:0] vwire_12_0;
	reg signed[17:0] vreg_12_0;
	node n12_0(.left(vreg_11_0), .right(vreg_13_0), .up(vreg_12_1), .down(vreg_12_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_0), .sw(sw));
	wire signed[17:0] vwire_12_1;
	reg signed[17:0] vreg_12_1;
	node n12_1(.left(vreg_11_1), .right(vreg_13_1), .up(vreg_12_2), .down(vreg_12_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_1), .sw(sw));
	wire signed[17:0] vwire_12_2;
	reg signed[17:0] vreg_12_2;
	node n12_2(.left(vreg_11_2), .right(vreg_13_2), .up(vreg_12_3), .down(vreg_12_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_2), .sw(sw));
	wire signed[17:0] vwire_12_3;
	reg signed[17:0] vreg_12_3;
	node n12_3(.left(vreg_11_3), .right(vreg_13_3), .up(vreg_12_4), .down(vreg_12_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_3), .sw(sw));
	wire signed[17:0] vwire_12_4;
	reg signed[17:0] vreg_12_4;
	node n12_4(.left(vreg_11_4), .right(vreg_13_4), .up(vreg_12_5), .down(vreg_12_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_4), .sw(sw));
	wire signed[17:0] vwire_12_5;
	reg signed[17:0] vreg_12_5;
	node n12_5(.left(vreg_11_5), .right(vreg_13_5), .up(vreg_12_6), .down(vreg_12_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_5), .sw(sw));
	wire signed[17:0] vwire_12_6;
	reg signed[17:0] vreg_12_6;
	node n12_6(.left(vreg_11_6), .right(vreg_13_6), .up(vreg_12_7), .down(vreg_12_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_6), .sw(sw));
	wire signed[17:0] vwire_12_7;
	reg signed[17:0] vreg_12_7;
	node n12_7(.left(vreg_11_7), .right(vreg_13_7), .up(vreg_12_8), .down(vreg_12_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_7), .sw(sw));
	wire signed[17:0] vwire_12_8;
	reg signed[17:0] vreg_12_8;
	node n12_8(.left(vreg_11_8), .right(vreg_13_8), .up(vreg_12_9), .down(vreg_12_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_8), .sw(sw));
	wire signed[17:0] vwire_12_9;
	reg signed[17:0] vreg_12_9;
	node n12_9(.left(vreg_11_9), .right(vreg_13_9), .up(vreg_12_10), .down(vreg_12_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_9), .sw(sw));
	wire signed[17:0] vwire_12_10;
	reg signed[17:0] vreg_12_10;
	node n12_10(.left(vreg_11_10), .right(vreg_13_10), .up(vreg_12_11), .down(vreg_12_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_10), .sw(sw));
	wire signed[17:0] vwire_12_11;
	reg signed[17:0] vreg_12_11;
	node n12_11(.left(vreg_11_11), .right(vreg_13_11), .up(vreg_12_12), .down(vreg_12_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_11), .sw(sw));
	wire signed[17:0] vwire_12_12;
	reg signed[17:0] vreg_12_12;
	node n12_12(.left(vreg_11_12), .right(vreg_13_12), .up(vreg_12_13), .down(vreg_12_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_12), .sw(sw));
	wire signed[17:0] vwire_12_13;
	reg signed[17:0] vreg_12_13;
	node n12_13(.left(vreg_11_13), .right(vreg_13_13), .up(vreg_12_14), .down(vreg_12_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_13), .sw(sw));
	wire signed[17:0] vwire_12_14;
	reg signed[17:0] vreg_12_14;
	node n12_14(.left(vreg_11_14), .right(vreg_13_14), .up(vreg_12_15), .down(vreg_12_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_14), .sw(sw));
	wire signed[17:0] vwire_12_15;
	reg signed[17:0] vreg_12_15;
	node n12_15(.left(vreg_11_15), .right(vreg_13_15), .up(vreg_12_16), .down(vreg_12_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_15), .sw(sw));
	wire signed[17:0] vwire_12_16;
	reg signed[17:0] vreg_12_16;
	node n12_16(.left(vreg_11_16), .right(vreg_13_16), .up(vreg_12_17), .down(vreg_12_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_16), .sw(sw));
	wire signed[17:0] vwire_12_17;
	reg signed[17:0] vreg_12_17;
	node n12_17(.left(vreg_11_17), .right(vreg_13_17), .up(vreg_12_18), .down(vreg_12_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_17), .sw(sw));
	wire signed[17:0] vwire_12_18;
	reg signed[17:0] vreg_12_18;
	node n12_18(.left(vreg_11_18), .right(vreg_13_18), .up(vreg_12_19), .down(vreg_12_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_18), .sw(sw));
	wire signed[17:0] vwire_12_19;
	reg signed[17:0] vreg_12_19;
	node n12_19(.left(vreg_11_19), .right(vreg_13_19), .up(vreg_12_20), .down(vreg_12_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_19), .sw(sw));
	wire signed[17:0] vwire_12_20;
	reg signed[17:0] vreg_12_20;
	node n12_20(.left(vreg_11_20), .right(vreg_13_20), .up(vreg_12_21), .down(vreg_12_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_20), .sw(sw));
	wire signed[17:0] vwire_12_21;
	reg signed[17:0] vreg_12_21;
	node n12_21(.left(vreg_11_21), .right(vreg_13_21), .up(vreg_12_22), .down(vreg_12_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_21), .sw(sw));
	wire signed[17:0] vwire_12_22;
	reg signed[17:0] vreg_12_22;
	node n12_22(.left(vreg_11_22), .right(vreg_13_22), .up(vreg_12_23), .down(vreg_12_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_22), .sw(sw));
	wire signed[17:0] vwire_12_23;
	reg signed[17:0] vreg_12_23;
	node n12_23(.left(vreg_11_23), .right(vreg_13_23), .up(vreg_12_24), .down(vreg_12_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_23), .sw(sw));
	wire signed[17:0] vwire_12_24;
	reg signed[17:0] vreg_12_24;
	node n12_24(.left(vreg_11_24), .right(vreg_13_24), .up(vreg_12_25), .down(vreg_12_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_24), .sw(sw));
	wire signed[17:0] vwire_12_25;
	reg signed[17:0] vreg_12_25;
	node n12_25(.left(vreg_11_25), .right(vreg_13_25), .up(vreg_12_26), .down(vreg_12_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_25), .sw(sw));
	wire signed[17:0] vwire_12_26;
	reg signed[17:0] vreg_12_26;
	node n12_26(.left(vreg_11_26), .right(vreg_13_26), .up(vreg_12_27), .down(vreg_12_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_26), .sw(sw));
	wire signed[17:0] vwire_12_27;
	reg signed[17:0] vreg_12_27;
	node n12_27(.left(vreg_11_27), .right(vreg_13_27), .up(vreg_12_28), .down(vreg_12_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_27), .sw(sw));
	wire signed[17:0] vwire_12_28;
	reg signed[17:0] vreg_12_28;
	node n12_28(.left(vreg_11_28), .right(vreg_13_28), .up(vreg_12_29), .down(vreg_12_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_28), .sw(sw));
	wire signed[17:0] vwire_12_29;
	reg signed[17:0] vreg_12_29;
	node n12_29(.left(vreg_11_29), .right(vreg_13_29), .up(vreg_12_30), .down(vreg_12_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_29), .sw(sw));
	wire signed[17:0] vwire_12_30;
	reg signed[17:0] vreg_12_30;
	node n12_30(.left(vreg_11_30), .right(vreg_13_30), .up(vreg_12_31), .down(vreg_12_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_30), .sw(sw));
	wire signed[17:0] vwire_12_31;
	reg signed[17:0] vreg_12_31;
	node n12_31(.left(vreg_11_31), .right(vreg_13_31), .up(vreg_12_32), .down(vreg_12_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_31), .sw(sw));
	wire signed[17:0] vwire_12_32;
	reg signed[17:0] vreg_12_32;
	node n12_32(.left(vreg_11_32), .right(vreg_13_32), .up(vreg_12_33), .down(vreg_12_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_32), .sw(sw));
	wire signed[17:0] vwire_12_33;
	reg signed[17:0] vreg_12_33;
	node n12_33(.left(vreg_11_33), .right(vreg_13_33), .up(vreg_12_34), .down(vreg_12_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_33), .sw(sw));
	wire signed[17:0] vwire_12_34;
	reg signed[17:0] vreg_12_34;
	node n12_34(.left(vreg_11_34), .right(vreg_13_34), .up(vreg_12_35), .down(vreg_12_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_34), .sw(sw));
	wire signed[17:0] vwire_12_35;
	reg signed[17:0] vreg_12_35;
	node n12_35(.left(vreg_11_35), .right(vreg_13_35), .up(vreg_12_36), .down(vreg_12_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_35), .sw(sw));
	wire signed[17:0] vwire_12_36;
	reg signed[17:0] vreg_12_36;
	node n12_36(.left(vreg_11_36), .right(vreg_13_36), .up(vreg_12_37), .down(vreg_12_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_36), .sw(sw));
	wire signed[17:0] vwire_12_37;
	reg signed[17:0] vreg_12_37;
	node n12_37(.left(vreg_11_37), .right(vreg_13_37), .up(vreg_12_38), .down(vreg_12_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_37), .sw(sw));
	wire signed[17:0] vwire_12_38;
	reg signed[17:0] vreg_12_38;
	node n12_38(.left(vreg_11_38), .right(vreg_13_38), .up(vreg_12_39), .down(vreg_12_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_38), .sw(sw));
	wire signed[17:0] vwire_12_39;
	reg signed[17:0] vreg_12_39;
	node n12_39(.left(vreg_11_39), .right(vreg_13_39), .up(vreg_12_40), .down(vreg_12_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_39), .sw(sw));
	wire signed[17:0] vwire_12_40;
	reg signed[17:0] vreg_12_40;
	node n12_40(.left(vreg_11_40), .right(vreg_13_40), .up(vreg_12_41), .down(vreg_12_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_40), .sw(sw));
	wire signed[17:0] vwire_12_41;
	reg signed[17:0] vreg_12_41;
	node n12_41(.left(vreg_11_41), .right(vreg_13_41), .up(vreg_12_42), .down(vreg_12_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_41), .sw(sw));
	wire signed[17:0] vwire_12_42;
	reg signed[17:0] vreg_12_42;
	node n12_42(.left(vreg_11_42), .right(vreg_13_42), .up(vreg_12_43), .down(vreg_12_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_42), .sw(sw));
	wire signed[17:0] vwire_12_43;
	reg signed[17:0] vreg_12_43;
	node n12_43(.left(vreg_11_43), .right(vreg_13_43), .up(vreg_12_44), .down(vreg_12_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_43), .sw(sw));
	wire signed[17:0] vwire_12_44;
	reg signed[17:0] vreg_12_44;
	node n12_44(.left(vreg_11_44), .right(vreg_13_44), .up(vreg_12_45), .down(vreg_12_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_44), .sw(sw));
	wire signed[17:0] vwire_12_45;
	reg signed[17:0] vreg_12_45;
	node n12_45(.left(vreg_11_45), .right(vreg_13_45), .up(vreg_12_46), .down(vreg_12_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_45), .sw(sw));
	wire signed[17:0] vwire_12_46;
	reg signed[17:0] vreg_12_46;
	node n12_46(.left(vreg_11_46), .right(vreg_13_46), .up(vreg_12_47), .down(vreg_12_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_46), .sw(sw));
	wire signed[17:0] vwire_12_47;
	reg signed[17:0] vreg_12_47;
	node n12_47(.left(vreg_11_47), .right(vreg_13_47), .up(vreg_12_48), .down(vreg_12_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_47), .sw(sw));
	wire signed[17:0] vwire_12_48;
	reg signed[17:0] vreg_12_48;
	node n12_48(.left(vreg_11_48), .right(vreg_13_48), .up(vreg_12_49), .down(vreg_12_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_48), .sw(sw));
	wire signed[17:0] vwire_12_49;
	reg signed[17:0] vreg_12_49;
	node n12_49(.left(vreg_11_49), .right(vreg_13_49), .up(18'b0), .down(vreg_12_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_12_49), .sw(sw));
	wire signed[17:0] vwire_13_0;
	reg signed[17:0] vreg_13_0;
	node n13_0(.left(vreg_12_0), .right(vreg_14_0), .up(vreg_13_1), .down(vreg_13_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_0), .sw(sw));
	wire signed[17:0] vwire_13_1;
	reg signed[17:0] vreg_13_1;
	node n13_1(.left(vreg_12_1), .right(vreg_14_1), .up(vreg_13_2), .down(vreg_13_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_1), .sw(sw));
	wire signed[17:0] vwire_13_2;
	reg signed[17:0] vreg_13_2;
	node n13_2(.left(vreg_12_2), .right(vreg_14_2), .up(vreg_13_3), .down(vreg_13_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_2), .sw(sw));
	wire signed[17:0] vwire_13_3;
	reg signed[17:0] vreg_13_3;
	node n13_3(.left(vreg_12_3), .right(vreg_14_3), .up(vreg_13_4), .down(vreg_13_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_3), .sw(sw));
	wire signed[17:0] vwire_13_4;
	reg signed[17:0] vreg_13_4;
	node n13_4(.left(vreg_12_4), .right(vreg_14_4), .up(vreg_13_5), .down(vreg_13_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_4), .sw(sw));
	wire signed[17:0] vwire_13_5;
	reg signed[17:0] vreg_13_5;
	node n13_5(.left(vreg_12_5), .right(vreg_14_5), .up(vreg_13_6), .down(vreg_13_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_5), .sw(sw));
	wire signed[17:0] vwire_13_6;
	reg signed[17:0] vreg_13_6;
	node n13_6(.left(vreg_12_6), .right(vreg_14_6), .up(vreg_13_7), .down(vreg_13_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_6), .sw(sw));
	wire signed[17:0] vwire_13_7;
	reg signed[17:0] vreg_13_7;
	node n13_7(.left(vreg_12_7), .right(vreg_14_7), .up(vreg_13_8), .down(vreg_13_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_7), .sw(sw));
	wire signed[17:0] vwire_13_8;
	reg signed[17:0] vreg_13_8;
	node n13_8(.left(vreg_12_8), .right(vreg_14_8), .up(vreg_13_9), .down(vreg_13_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_8), .sw(sw));
	wire signed[17:0] vwire_13_9;
	reg signed[17:0] vreg_13_9;
	node n13_9(.left(vreg_12_9), .right(vreg_14_9), .up(vreg_13_10), .down(vreg_13_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_9), .sw(sw));
	wire signed[17:0] vwire_13_10;
	reg signed[17:0] vreg_13_10;
	node n13_10(.left(vreg_12_10), .right(vreg_14_10), .up(vreg_13_11), .down(vreg_13_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_10), .sw(sw));
	wire signed[17:0] vwire_13_11;
	reg signed[17:0] vreg_13_11;
	node n13_11(.left(vreg_12_11), .right(vreg_14_11), .up(vreg_13_12), .down(vreg_13_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_11), .sw(sw));
	wire signed[17:0] vwire_13_12;
	reg signed[17:0] vreg_13_12;
	node n13_12(.left(vreg_12_12), .right(vreg_14_12), .up(vreg_13_13), .down(vreg_13_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_12), .sw(sw));
	wire signed[17:0] vwire_13_13;
	reg signed[17:0] vreg_13_13;
	node n13_13(.left(vreg_12_13), .right(vreg_14_13), .up(vreg_13_14), .down(vreg_13_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_13), .sw(sw));
	wire signed[17:0] vwire_13_14;
	reg signed[17:0] vreg_13_14;
	node n13_14(.left(vreg_12_14), .right(vreg_14_14), .up(vreg_13_15), .down(vreg_13_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_14), .sw(sw));
	wire signed[17:0] vwire_13_15;
	reg signed[17:0] vreg_13_15;
	node n13_15(.left(vreg_12_15), .right(vreg_14_15), .up(vreg_13_16), .down(vreg_13_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_15), .sw(sw));
	wire signed[17:0] vwire_13_16;
	reg signed[17:0] vreg_13_16;
	node n13_16(.left(vreg_12_16), .right(vreg_14_16), .up(vreg_13_17), .down(vreg_13_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_16), .sw(sw));
	wire signed[17:0] vwire_13_17;
	reg signed[17:0] vreg_13_17;
	node n13_17(.left(vreg_12_17), .right(vreg_14_17), .up(vreg_13_18), .down(vreg_13_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_17), .sw(sw));
	wire signed[17:0] vwire_13_18;
	reg signed[17:0] vreg_13_18;
	node n13_18(.left(vreg_12_18), .right(vreg_14_18), .up(vreg_13_19), .down(vreg_13_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_18), .sw(sw));
	wire signed[17:0] vwire_13_19;
	reg signed[17:0] vreg_13_19;
	node n13_19(.left(vreg_12_19), .right(vreg_14_19), .up(vreg_13_20), .down(vreg_13_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_19), .sw(sw));
	wire signed[17:0] vwire_13_20;
	reg signed[17:0] vreg_13_20;
	node n13_20(.left(vreg_12_20), .right(vreg_14_20), .up(vreg_13_21), .down(vreg_13_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_20), .sw(sw));
	wire signed[17:0] vwire_13_21;
	reg signed[17:0] vreg_13_21;
	node n13_21(.left(vreg_12_21), .right(vreg_14_21), .up(vreg_13_22), .down(vreg_13_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_21), .sw(sw));
	wire signed[17:0] vwire_13_22;
	reg signed[17:0] vreg_13_22;
	node n13_22(.left(vreg_12_22), .right(vreg_14_22), .up(vreg_13_23), .down(vreg_13_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_22), .sw(sw));
	wire signed[17:0] vwire_13_23;
	reg signed[17:0] vreg_13_23;
	node n13_23(.left(vreg_12_23), .right(vreg_14_23), .up(vreg_13_24), .down(vreg_13_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_23), .sw(sw));
	wire signed[17:0] vwire_13_24;
	reg signed[17:0] vreg_13_24;
	node n13_24(.left(vreg_12_24), .right(vreg_14_24), .up(vreg_13_25), .down(vreg_13_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_24), .sw(sw));
	wire signed[17:0] vwire_13_25;
	reg signed[17:0] vreg_13_25;
	node n13_25(.left(vreg_12_25), .right(vreg_14_25), .up(vreg_13_26), .down(vreg_13_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_25), .sw(sw));
	wire signed[17:0] vwire_13_26;
	reg signed[17:0] vreg_13_26;
	node n13_26(.left(vreg_12_26), .right(vreg_14_26), .up(vreg_13_27), .down(vreg_13_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_26), .sw(sw));
	wire signed[17:0] vwire_13_27;
	reg signed[17:0] vreg_13_27;
	node n13_27(.left(vreg_12_27), .right(vreg_14_27), .up(vreg_13_28), .down(vreg_13_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_27), .sw(sw));
	wire signed[17:0] vwire_13_28;
	reg signed[17:0] vreg_13_28;
	node n13_28(.left(vreg_12_28), .right(vreg_14_28), .up(vreg_13_29), .down(vreg_13_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_28), .sw(sw));
	wire signed[17:0] vwire_13_29;
	reg signed[17:0] vreg_13_29;
	node n13_29(.left(vreg_12_29), .right(vreg_14_29), .up(vreg_13_30), .down(vreg_13_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_29), .sw(sw));
	wire signed[17:0] vwire_13_30;
	reg signed[17:0] vreg_13_30;
	node n13_30(.left(vreg_12_30), .right(vreg_14_30), .up(vreg_13_31), .down(vreg_13_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_30), .sw(sw));
	wire signed[17:0] vwire_13_31;
	reg signed[17:0] vreg_13_31;
	node n13_31(.left(vreg_12_31), .right(vreg_14_31), .up(vreg_13_32), .down(vreg_13_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_31), .sw(sw));
	wire signed[17:0] vwire_13_32;
	reg signed[17:0] vreg_13_32;
	node n13_32(.left(vreg_12_32), .right(vreg_14_32), .up(vreg_13_33), .down(vreg_13_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_32), .sw(sw));
	wire signed[17:0] vwire_13_33;
	reg signed[17:0] vreg_13_33;
	node n13_33(.left(vreg_12_33), .right(vreg_14_33), .up(vreg_13_34), .down(vreg_13_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_33), .sw(sw));
	wire signed[17:0] vwire_13_34;
	reg signed[17:0] vreg_13_34;
	node n13_34(.left(vreg_12_34), .right(vreg_14_34), .up(vreg_13_35), .down(vreg_13_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_34), .sw(sw));
	wire signed[17:0] vwire_13_35;
	reg signed[17:0] vreg_13_35;
	node n13_35(.left(vreg_12_35), .right(vreg_14_35), .up(vreg_13_36), .down(vreg_13_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_35), .sw(sw));
	wire signed[17:0] vwire_13_36;
	reg signed[17:0] vreg_13_36;
	node n13_36(.left(vreg_12_36), .right(vreg_14_36), .up(vreg_13_37), .down(vreg_13_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_36), .sw(sw));
	wire signed[17:0] vwire_13_37;
	reg signed[17:0] vreg_13_37;
	node n13_37(.left(vreg_12_37), .right(vreg_14_37), .up(vreg_13_38), .down(vreg_13_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_37), .sw(sw));
	wire signed[17:0] vwire_13_38;
	reg signed[17:0] vreg_13_38;
	node n13_38(.left(vreg_12_38), .right(vreg_14_38), .up(vreg_13_39), .down(vreg_13_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_38), .sw(sw));
	wire signed[17:0] vwire_13_39;
	reg signed[17:0] vreg_13_39;
	node n13_39(.left(vreg_12_39), .right(vreg_14_39), .up(vreg_13_40), .down(vreg_13_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_39), .sw(sw));
	wire signed[17:0] vwire_13_40;
	reg signed[17:0] vreg_13_40;
	node n13_40(.left(vreg_12_40), .right(vreg_14_40), .up(vreg_13_41), .down(vreg_13_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_40), .sw(sw));
	wire signed[17:0] vwire_13_41;
	reg signed[17:0] vreg_13_41;
	node n13_41(.left(vreg_12_41), .right(vreg_14_41), .up(vreg_13_42), .down(vreg_13_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_41), .sw(sw));
	wire signed[17:0] vwire_13_42;
	reg signed[17:0] vreg_13_42;
	node n13_42(.left(vreg_12_42), .right(vreg_14_42), .up(vreg_13_43), .down(vreg_13_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_42), .sw(sw));
	wire signed[17:0] vwire_13_43;
	reg signed[17:0] vreg_13_43;
	node n13_43(.left(vreg_12_43), .right(vreg_14_43), .up(vreg_13_44), .down(vreg_13_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_43), .sw(sw));
	wire signed[17:0] vwire_13_44;
	reg signed[17:0] vreg_13_44;
	node n13_44(.left(vreg_12_44), .right(vreg_14_44), .up(vreg_13_45), .down(vreg_13_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_44), .sw(sw));
	wire signed[17:0] vwire_13_45;
	reg signed[17:0] vreg_13_45;
	node n13_45(.left(vreg_12_45), .right(vreg_14_45), .up(vreg_13_46), .down(vreg_13_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_45), .sw(sw));
	wire signed[17:0] vwire_13_46;
	reg signed[17:0] vreg_13_46;
	node n13_46(.left(vreg_12_46), .right(vreg_14_46), .up(vreg_13_47), .down(vreg_13_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_46), .sw(sw));
	wire signed[17:0] vwire_13_47;
	reg signed[17:0] vreg_13_47;
	node n13_47(.left(vreg_12_47), .right(vreg_14_47), .up(vreg_13_48), .down(vreg_13_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_47), .sw(sw));
	wire signed[17:0] vwire_13_48;
	reg signed[17:0] vreg_13_48;
	node n13_48(.left(vreg_12_48), .right(vreg_14_48), .up(vreg_13_49), .down(vreg_13_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_48), .sw(sw));
	wire signed[17:0] vwire_13_49;
	reg signed[17:0] vreg_13_49;
	node n13_49(.left(vreg_12_49), .right(vreg_14_49), .up(18'b0), .down(vreg_13_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_13_49), .sw(sw));
	wire signed[17:0] vwire_14_0;
	reg signed[17:0] vreg_14_0;
	node n14_0(.left(vreg_13_0), .right(vreg_15_0), .up(vreg_14_1), .down(vreg_14_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_0), .sw(sw));
	wire signed[17:0] vwire_14_1;
	reg signed[17:0] vreg_14_1;
	node n14_1(.left(vreg_13_1), .right(vreg_15_1), .up(vreg_14_2), .down(vreg_14_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_1), .sw(sw));
	wire signed[17:0] vwire_14_2;
	reg signed[17:0] vreg_14_2;
	node n14_2(.left(vreg_13_2), .right(vreg_15_2), .up(vreg_14_3), .down(vreg_14_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_2), .sw(sw));
	wire signed[17:0] vwire_14_3;
	reg signed[17:0] vreg_14_3;
	node n14_3(.left(vreg_13_3), .right(vreg_15_3), .up(vreg_14_4), .down(vreg_14_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_3), .sw(sw));
	wire signed[17:0] vwire_14_4;
	reg signed[17:0] vreg_14_4;
	node n14_4(.left(vreg_13_4), .right(vreg_15_4), .up(vreg_14_5), .down(vreg_14_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_4), .sw(sw));
	wire signed[17:0] vwire_14_5;
	reg signed[17:0] vreg_14_5;
	node n14_5(.left(vreg_13_5), .right(vreg_15_5), .up(vreg_14_6), .down(vreg_14_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_5), .sw(sw));
	wire signed[17:0] vwire_14_6;
	reg signed[17:0] vreg_14_6;
	node n14_6(.left(vreg_13_6), .right(vreg_15_6), .up(vreg_14_7), .down(vreg_14_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_6), .sw(sw));
	wire signed[17:0] vwire_14_7;
	reg signed[17:0] vreg_14_7;
	node n14_7(.left(vreg_13_7), .right(vreg_15_7), .up(vreg_14_8), .down(vreg_14_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_7), .sw(sw));
	wire signed[17:0] vwire_14_8;
	reg signed[17:0] vreg_14_8;
	node n14_8(.left(vreg_13_8), .right(vreg_15_8), .up(vreg_14_9), .down(vreg_14_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_8), .sw(sw));
	wire signed[17:0] vwire_14_9;
	reg signed[17:0] vreg_14_9;
	node n14_9(.left(vreg_13_9), .right(vreg_15_9), .up(vreg_14_10), .down(vreg_14_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_9), .sw(sw));
	wire signed[17:0] vwire_14_10;
	reg signed[17:0] vreg_14_10;
	node n14_10(.left(vreg_13_10), .right(vreg_15_10), .up(vreg_14_11), .down(vreg_14_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_10), .sw(sw));
	wire signed[17:0] vwire_14_11;
	reg signed[17:0] vreg_14_11;
	node n14_11(.left(vreg_13_11), .right(vreg_15_11), .up(vreg_14_12), .down(vreg_14_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_11), .sw(sw));
	wire signed[17:0] vwire_14_12;
	reg signed[17:0] vreg_14_12;
	node n14_12(.left(vreg_13_12), .right(vreg_15_12), .up(vreg_14_13), .down(vreg_14_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_12), .sw(sw));
	wire signed[17:0] vwire_14_13;
	reg signed[17:0] vreg_14_13;
	node n14_13(.left(vreg_13_13), .right(vreg_15_13), .up(vreg_14_14), .down(vreg_14_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_13), .sw(sw));
	wire signed[17:0] vwire_14_14;
	reg signed[17:0] vreg_14_14;
	node n14_14(.left(vreg_13_14), .right(vreg_15_14), .up(vreg_14_15), .down(vreg_14_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_14), .sw(sw));
	wire signed[17:0] vwire_14_15;
	reg signed[17:0] vreg_14_15;
	node n14_15(.left(vreg_13_15), .right(vreg_15_15), .up(vreg_14_16), .down(vreg_14_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_15), .sw(sw));
	wire signed[17:0] vwire_14_16;
	reg signed[17:0] vreg_14_16;
	node n14_16(.left(vreg_13_16), .right(vreg_15_16), .up(vreg_14_17), .down(vreg_14_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_16), .sw(sw));
	wire signed[17:0] vwire_14_17;
	reg signed[17:0] vreg_14_17;
	node n14_17(.left(vreg_13_17), .right(vreg_15_17), .up(vreg_14_18), .down(vreg_14_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_17), .sw(sw));
	wire signed[17:0] vwire_14_18;
	reg signed[17:0] vreg_14_18;
	node n14_18(.left(vreg_13_18), .right(vreg_15_18), .up(vreg_14_19), .down(vreg_14_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_18), .sw(sw));
	wire signed[17:0] vwire_14_19;
	reg signed[17:0] vreg_14_19;
	node n14_19(.left(vreg_13_19), .right(vreg_15_19), .up(vreg_14_20), .down(vreg_14_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_19), .sw(sw));
	wire signed[17:0] vwire_14_20;
	reg signed[17:0] vreg_14_20;
	node n14_20(.left(vreg_13_20), .right(vreg_15_20), .up(vreg_14_21), .down(vreg_14_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_20), .sw(sw));
	wire signed[17:0] vwire_14_21;
	reg signed[17:0] vreg_14_21;
	node n14_21(.left(vreg_13_21), .right(vreg_15_21), .up(vreg_14_22), .down(vreg_14_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_21), .sw(sw));
	wire signed[17:0] vwire_14_22;
	reg signed[17:0] vreg_14_22;
	node n14_22(.left(vreg_13_22), .right(vreg_15_22), .up(vreg_14_23), .down(vreg_14_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_22), .sw(sw));
	wire signed[17:0] vwire_14_23;
	reg signed[17:0] vreg_14_23;
	node n14_23(.left(vreg_13_23), .right(vreg_15_23), .up(vreg_14_24), .down(vreg_14_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_23), .sw(sw));
	wire signed[17:0] vwire_14_24;
	reg signed[17:0] vreg_14_24;
	node n14_24(.left(vreg_13_24), .right(vreg_15_24), .up(vreg_14_25), .down(vreg_14_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_24), .sw(sw));
	wire signed[17:0] vwire_14_25;
	reg signed[17:0] vreg_14_25;
	node n14_25(.left(vreg_13_25), .right(vreg_15_25), .up(vreg_14_26), .down(vreg_14_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_25), .sw(sw));
	wire signed[17:0] vwire_14_26;
	reg signed[17:0] vreg_14_26;
	node n14_26(.left(vreg_13_26), .right(vreg_15_26), .up(vreg_14_27), .down(vreg_14_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_26), .sw(sw));
	wire signed[17:0] vwire_14_27;
	reg signed[17:0] vreg_14_27;
	node n14_27(.left(vreg_13_27), .right(vreg_15_27), .up(vreg_14_28), .down(vreg_14_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_27), .sw(sw));
	wire signed[17:0] vwire_14_28;
	reg signed[17:0] vreg_14_28;
	node n14_28(.left(vreg_13_28), .right(vreg_15_28), .up(vreg_14_29), .down(vreg_14_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_28), .sw(sw));
	wire signed[17:0] vwire_14_29;
	reg signed[17:0] vreg_14_29;
	node n14_29(.left(vreg_13_29), .right(vreg_15_29), .up(vreg_14_30), .down(vreg_14_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_29), .sw(sw));
	wire signed[17:0] vwire_14_30;
	reg signed[17:0] vreg_14_30;
	node n14_30(.left(vreg_13_30), .right(vreg_15_30), .up(vreg_14_31), .down(vreg_14_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_30), .sw(sw));
	wire signed[17:0] vwire_14_31;
	reg signed[17:0] vreg_14_31;
	node n14_31(.left(vreg_13_31), .right(vreg_15_31), .up(vreg_14_32), .down(vreg_14_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_31), .sw(sw));
	wire signed[17:0] vwire_14_32;
	reg signed[17:0] vreg_14_32;
	node n14_32(.left(vreg_13_32), .right(vreg_15_32), .up(vreg_14_33), .down(vreg_14_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_32), .sw(sw));
	wire signed[17:0] vwire_14_33;
	reg signed[17:0] vreg_14_33;
	node n14_33(.left(vreg_13_33), .right(vreg_15_33), .up(vreg_14_34), .down(vreg_14_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_33), .sw(sw));
	wire signed[17:0] vwire_14_34;
	reg signed[17:0] vreg_14_34;
	node n14_34(.left(vreg_13_34), .right(vreg_15_34), .up(vreg_14_35), .down(vreg_14_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_34), .sw(sw));
	wire signed[17:0] vwire_14_35;
	reg signed[17:0] vreg_14_35;
	node n14_35(.left(vreg_13_35), .right(vreg_15_35), .up(vreg_14_36), .down(vreg_14_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_35), .sw(sw));
	wire signed[17:0] vwire_14_36;
	reg signed[17:0] vreg_14_36;
	node n14_36(.left(vreg_13_36), .right(vreg_15_36), .up(vreg_14_37), .down(vreg_14_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_36), .sw(sw));
	wire signed[17:0] vwire_14_37;
	reg signed[17:0] vreg_14_37;
	node n14_37(.left(vreg_13_37), .right(vreg_15_37), .up(vreg_14_38), .down(vreg_14_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_37), .sw(sw));
	wire signed[17:0] vwire_14_38;
	reg signed[17:0] vreg_14_38;
	node n14_38(.left(vreg_13_38), .right(vreg_15_38), .up(vreg_14_39), .down(vreg_14_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_38), .sw(sw));
	wire signed[17:0] vwire_14_39;
	reg signed[17:0] vreg_14_39;
	node n14_39(.left(vreg_13_39), .right(vreg_15_39), .up(vreg_14_40), .down(vreg_14_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_39), .sw(sw));
	wire signed[17:0] vwire_14_40;
	reg signed[17:0] vreg_14_40;
	node n14_40(.left(vreg_13_40), .right(vreg_15_40), .up(vreg_14_41), .down(vreg_14_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_40), .sw(sw));
	wire signed[17:0] vwire_14_41;
	reg signed[17:0] vreg_14_41;
	node n14_41(.left(vreg_13_41), .right(vreg_15_41), .up(vreg_14_42), .down(vreg_14_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_41), .sw(sw));
	wire signed[17:0] vwire_14_42;
	reg signed[17:0] vreg_14_42;
	node n14_42(.left(vreg_13_42), .right(vreg_15_42), .up(vreg_14_43), .down(vreg_14_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_42), .sw(sw));
	wire signed[17:0] vwire_14_43;
	reg signed[17:0] vreg_14_43;
	node n14_43(.left(vreg_13_43), .right(vreg_15_43), .up(vreg_14_44), .down(vreg_14_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_43), .sw(sw));
	wire signed[17:0] vwire_14_44;
	reg signed[17:0] vreg_14_44;
	node n14_44(.left(vreg_13_44), .right(vreg_15_44), .up(vreg_14_45), .down(vreg_14_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_44), .sw(sw));
	wire signed[17:0] vwire_14_45;
	reg signed[17:0] vreg_14_45;
	node n14_45(.left(vreg_13_45), .right(vreg_15_45), .up(vreg_14_46), .down(vreg_14_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_45), .sw(sw));
	wire signed[17:0] vwire_14_46;
	reg signed[17:0] vreg_14_46;
	node n14_46(.left(vreg_13_46), .right(vreg_15_46), .up(vreg_14_47), .down(vreg_14_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_46), .sw(sw));
	wire signed[17:0] vwire_14_47;
	reg signed[17:0] vreg_14_47;
	node n14_47(.left(vreg_13_47), .right(vreg_15_47), .up(vreg_14_48), .down(vreg_14_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_47), .sw(sw));
	wire signed[17:0] vwire_14_48;
	reg signed[17:0] vreg_14_48;
	node n14_48(.left(vreg_13_48), .right(vreg_15_48), .up(vreg_14_49), .down(vreg_14_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_48), .sw(sw));
	wire signed[17:0] vwire_14_49;
	reg signed[17:0] vreg_14_49;
	node n14_49(.left(vreg_13_49), .right(vreg_15_49), .up(18'b0), .down(vreg_14_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_14_49), .sw(sw));
	wire signed[17:0] vwire_15_0;
	reg signed[17:0] vreg_15_0;
	node n15_0(.left(vreg_14_0), .right(vreg_16_0), .up(vreg_15_1), .down(vreg_15_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_0), .sw(sw));
	wire signed[17:0] vwire_15_1;
	reg signed[17:0] vreg_15_1;
	node n15_1(.left(vreg_14_1), .right(vreg_16_1), .up(vreg_15_2), .down(vreg_15_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_1), .sw(sw));
	wire signed[17:0] vwire_15_2;
	reg signed[17:0] vreg_15_2;
	node n15_2(.left(vreg_14_2), .right(vreg_16_2), .up(vreg_15_3), .down(vreg_15_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_2), .sw(sw));
	wire signed[17:0] vwire_15_3;
	reg signed[17:0] vreg_15_3;
	node n15_3(.left(vreg_14_3), .right(vreg_16_3), .up(vreg_15_4), .down(vreg_15_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_3), .sw(sw));
	wire signed[17:0] vwire_15_4;
	reg signed[17:0] vreg_15_4;
	node n15_4(.left(vreg_14_4), .right(vreg_16_4), .up(vreg_15_5), .down(vreg_15_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_4), .sw(sw));
	wire signed[17:0] vwire_15_5;
	reg signed[17:0] vreg_15_5;
	node n15_5(.left(vreg_14_5), .right(vreg_16_5), .up(vreg_15_6), .down(vreg_15_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_5), .sw(sw));
	wire signed[17:0] vwire_15_6;
	reg signed[17:0] vreg_15_6;
	node n15_6(.left(vreg_14_6), .right(vreg_16_6), .up(vreg_15_7), .down(vreg_15_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_6), .sw(sw));
	wire signed[17:0] vwire_15_7;
	reg signed[17:0] vreg_15_7;
	node n15_7(.left(vreg_14_7), .right(vreg_16_7), .up(vreg_15_8), .down(vreg_15_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_7), .sw(sw));
	wire signed[17:0] vwire_15_8;
	reg signed[17:0] vreg_15_8;
	node n15_8(.left(vreg_14_8), .right(vreg_16_8), .up(vreg_15_9), .down(vreg_15_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_8), .sw(sw));
	wire signed[17:0] vwire_15_9;
	reg signed[17:0] vreg_15_9;
	node n15_9(.left(vreg_14_9), .right(vreg_16_9), .up(vreg_15_10), .down(vreg_15_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_9), .sw(sw));
	wire signed[17:0] vwire_15_10;
	reg signed[17:0] vreg_15_10;
	node n15_10(.left(vreg_14_10), .right(vreg_16_10), .up(vreg_15_11), .down(vreg_15_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_10), .sw(sw));
	wire signed[17:0] vwire_15_11;
	reg signed[17:0] vreg_15_11;
	node n15_11(.left(vreg_14_11), .right(vreg_16_11), .up(vreg_15_12), .down(vreg_15_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_11), .sw(sw));
	wire signed[17:0] vwire_15_12;
	reg signed[17:0] vreg_15_12;
	node n15_12(.left(vreg_14_12), .right(vreg_16_12), .up(vreg_15_13), .down(vreg_15_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_12), .sw(sw));
	wire signed[17:0] vwire_15_13;
	reg signed[17:0] vreg_15_13;
	node n15_13(.left(vreg_14_13), .right(vreg_16_13), .up(vreg_15_14), .down(vreg_15_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_13), .sw(sw));
	wire signed[17:0] vwire_15_14;
	reg signed[17:0] vreg_15_14;
	node n15_14(.left(vreg_14_14), .right(vreg_16_14), .up(vreg_15_15), .down(vreg_15_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_14), .sw(sw));
	wire signed[17:0] vwire_15_15;
	reg signed[17:0] vreg_15_15;
	node n15_15(.left(vreg_14_15), .right(vreg_16_15), .up(vreg_15_16), .down(vreg_15_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_15), .sw(sw));
	wire signed[17:0] vwire_15_16;
	reg signed[17:0] vreg_15_16;
	node n15_16(.left(vreg_14_16), .right(vreg_16_16), .up(vreg_15_17), .down(vreg_15_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_16), .sw(sw));
	wire signed[17:0] vwire_15_17;
	reg signed[17:0] vreg_15_17;
	node n15_17(.left(vreg_14_17), .right(vreg_16_17), .up(vreg_15_18), .down(vreg_15_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_17), .sw(sw));
	wire signed[17:0] vwire_15_18;
	reg signed[17:0] vreg_15_18;
	node n15_18(.left(vreg_14_18), .right(vreg_16_18), .up(vreg_15_19), .down(vreg_15_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_18), .sw(sw));
	wire signed[17:0] vwire_15_19;
	reg signed[17:0] vreg_15_19;
	node n15_19(.left(vreg_14_19), .right(vreg_16_19), .up(vreg_15_20), .down(vreg_15_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_19), .sw(sw));
	wire signed[17:0] vwire_15_20;
	reg signed[17:0] vreg_15_20;
	node n15_20(.left(vreg_14_20), .right(vreg_16_20), .up(vreg_15_21), .down(vreg_15_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_20), .sw(sw));
	wire signed[17:0] vwire_15_21;
	reg signed[17:0] vreg_15_21;
	node n15_21(.left(vreg_14_21), .right(vreg_16_21), .up(vreg_15_22), .down(vreg_15_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_21), .sw(sw));
	wire signed[17:0] vwire_15_22;
	reg signed[17:0] vreg_15_22;
	node n15_22(.left(vreg_14_22), .right(vreg_16_22), .up(vreg_15_23), .down(vreg_15_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_22), .sw(sw));
	wire signed[17:0] vwire_15_23;
	reg signed[17:0] vreg_15_23;
	node n15_23(.left(vreg_14_23), .right(vreg_16_23), .up(vreg_15_24), .down(vreg_15_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_23), .sw(sw));
	wire signed[17:0] vwire_15_24;
	reg signed[17:0] vreg_15_24;
	node n15_24(.left(vreg_14_24), .right(vreg_16_24), .up(vreg_15_25), .down(vreg_15_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_24), .sw(sw));
	wire signed[17:0] vwire_15_25;
	reg signed[17:0] vreg_15_25;
	node n15_25(.left(vreg_14_25), .right(vreg_16_25), .up(vreg_15_26), .down(vreg_15_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_25), .sw(sw));
	wire signed[17:0] vwire_15_26;
	reg signed[17:0] vreg_15_26;
	node n15_26(.left(vreg_14_26), .right(vreg_16_26), .up(vreg_15_27), .down(vreg_15_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_26), .sw(sw));
	wire signed[17:0] vwire_15_27;
	reg signed[17:0] vreg_15_27;
	node n15_27(.left(vreg_14_27), .right(vreg_16_27), .up(vreg_15_28), .down(vreg_15_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_27), .sw(sw));
	wire signed[17:0] vwire_15_28;
	reg signed[17:0] vreg_15_28;
	node n15_28(.left(vreg_14_28), .right(vreg_16_28), .up(vreg_15_29), .down(vreg_15_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_28), .sw(sw));
	wire signed[17:0] vwire_15_29;
	reg signed[17:0] vreg_15_29;
	node n15_29(.left(vreg_14_29), .right(vreg_16_29), .up(vreg_15_30), .down(vreg_15_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_29), .sw(sw));
	wire signed[17:0] vwire_15_30;
	reg signed[17:0] vreg_15_30;
	node n15_30(.left(vreg_14_30), .right(vreg_16_30), .up(vreg_15_31), .down(vreg_15_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_30), .sw(sw));
	wire signed[17:0] vwire_15_31;
	reg signed[17:0] vreg_15_31;
	node n15_31(.left(vreg_14_31), .right(vreg_16_31), .up(vreg_15_32), .down(vreg_15_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_31), .sw(sw));
	wire signed[17:0] vwire_15_32;
	reg signed[17:0] vreg_15_32;
	node n15_32(.left(vreg_14_32), .right(vreg_16_32), .up(vreg_15_33), .down(vreg_15_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_32), .sw(sw));
	wire signed[17:0] vwire_15_33;
	reg signed[17:0] vreg_15_33;
	node n15_33(.left(vreg_14_33), .right(vreg_16_33), .up(vreg_15_34), .down(vreg_15_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_33), .sw(sw));
	wire signed[17:0] vwire_15_34;
	reg signed[17:0] vreg_15_34;
	node n15_34(.left(vreg_14_34), .right(vreg_16_34), .up(vreg_15_35), .down(vreg_15_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_34), .sw(sw));
	wire signed[17:0] vwire_15_35;
	reg signed[17:0] vreg_15_35;
	node n15_35(.left(vreg_14_35), .right(vreg_16_35), .up(vreg_15_36), .down(vreg_15_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_35), .sw(sw));
	wire signed[17:0] vwire_15_36;
	reg signed[17:0] vreg_15_36;
	node n15_36(.left(vreg_14_36), .right(vreg_16_36), .up(vreg_15_37), .down(vreg_15_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_36), .sw(sw));
	wire signed[17:0] vwire_15_37;
	reg signed[17:0] vreg_15_37;
	node n15_37(.left(vreg_14_37), .right(vreg_16_37), .up(vreg_15_38), .down(vreg_15_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_37), .sw(sw));
	wire signed[17:0] vwire_15_38;
	reg signed[17:0] vreg_15_38;
	node n15_38(.left(vreg_14_38), .right(vreg_16_38), .up(vreg_15_39), .down(vreg_15_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_38), .sw(sw));
	wire signed[17:0] vwire_15_39;
	reg signed[17:0] vreg_15_39;
	node n15_39(.left(vreg_14_39), .right(vreg_16_39), .up(vreg_15_40), .down(vreg_15_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_39), .sw(sw));
	wire signed[17:0] vwire_15_40;
	reg signed[17:0] vreg_15_40;
	node n15_40(.left(vreg_14_40), .right(vreg_16_40), .up(vreg_15_41), .down(vreg_15_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_40), .sw(sw));
	wire signed[17:0] vwire_15_41;
	reg signed[17:0] vreg_15_41;
	node n15_41(.left(vreg_14_41), .right(vreg_16_41), .up(vreg_15_42), .down(vreg_15_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_41), .sw(sw));
	wire signed[17:0] vwire_15_42;
	reg signed[17:0] vreg_15_42;
	node n15_42(.left(vreg_14_42), .right(vreg_16_42), .up(vreg_15_43), .down(vreg_15_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_42), .sw(sw));
	wire signed[17:0] vwire_15_43;
	reg signed[17:0] vreg_15_43;
	node n15_43(.left(vreg_14_43), .right(vreg_16_43), .up(vreg_15_44), .down(vreg_15_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_43), .sw(sw));
	wire signed[17:0] vwire_15_44;
	reg signed[17:0] vreg_15_44;
	node n15_44(.left(vreg_14_44), .right(vreg_16_44), .up(vreg_15_45), .down(vreg_15_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_44), .sw(sw));
	wire signed[17:0] vwire_15_45;
	reg signed[17:0] vreg_15_45;
	node n15_45(.left(vreg_14_45), .right(vreg_16_45), .up(vreg_15_46), .down(vreg_15_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_45), .sw(sw));
	wire signed[17:0] vwire_15_46;
	reg signed[17:0] vreg_15_46;
	node n15_46(.left(vreg_14_46), .right(vreg_16_46), .up(vreg_15_47), .down(vreg_15_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_46), .sw(sw));
	wire signed[17:0] vwire_15_47;
	reg signed[17:0] vreg_15_47;
	node n15_47(.left(vreg_14_47), .right(vreg_16_47), .up(vreg_15_48), .down(vreg_15_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_47), .sw(sw));
	wire signed[17:0] vwire_15_48;
	reg signed[17:0] vreg_15_48;
	node n15_48(.left(vreg_14_48), .right(vreg_16_48), .up(vreg_15_49), .down(vreg_15_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_48), .sw(sw));
	wire signed[17:0] vwire_15_49;
	reg signed[17:0] vreg_15_49;
	node n15_49(.left(vreg_14_49), .right(vreg_16_49), .up(18'b0), .down(vreg_15_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_15_49), .sw(sw));
	wire signed[17:0] vwire_16_0;
	reg signed[17:0] vreg_16_0;
	node n16_0(.left(vreg_15_0), .right(vreg_17_0), .up(vreg_16_1), .down(vreg_16_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_0), .sw(sw));
	wire signed[17:0] vwire_16_1;
	reg signed[17:0] vreg_16_1;
	node n16_1(.left(vreg_15_1), .right(vreg_17_1), .up(vreg_16_2), .down(vreg_16_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_1), .sw(sw));
	wire signed[17:0] vwire_16_2;
	reg signed[17:0] vreg_16_2;
	node n16_2(.left(vreg_15_2), .right(vreg_17_2), .up(vreg_16_3), .down(vreg_16_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_2), .sw(sw));
	wire signed[17:0] vwire_16_3;
	reg signed[17:0] vreg_16_3;
	node n16_3(.left(vreg_15_3), .right(vreg_17_3), .up(vreg_16_4), .down(vreg_16_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_3), .sw(sw));
	wire signed[17:0] vwire_16_4;
	reg signed[17:0] vreg_16_4;
	node n16_4(.left(vreg_15_4), .right(vreg_17_4), .up(vreg_16_5), .down(vreg_16_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_4), .sw(sw));
	wire signed[17:0] vwire_16_5;
	reg signed[17:0] vreg_16_5;
	node n16_5(.left(vreg_15_5), .right(vreg_17_5), .up(vreg_16_6), .down(vreg_16_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_5), .sw(sw));
	wire signed[17:0] vwire_16_6;
	reg signed[17:0] vreg_16_6;
	node n16_6(.left(vreg_15_6), .right(vreg_17_6), .up(vreg_16_7), .down(vreg_16_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_6), .sw(sw));
	wire signed[17:0] vwire_16_7;
	reg signed[17:0] vreg_16_7;
	node n16_7(.left(vreg_15_7), .right(vreg_17_7), .up(vreg_16_8), .down(vreg_16_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_7), .sw(sw));
	wire signed[17:0] vwire_16_8;
	reg signed[17:0] vreg_16_8;
	node n16_8(.left(vreg_15_8), .right(vreg_17_8), .up(vreg_16_9), .down(vreg_16_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_8), .sw(sw));
	wire signed[17:0] vwire_16_9;
	reg signed[17:0] vreg_16_9;
	node n16_9(.left(vreg_15_9), .right(vreg_17_9), .up(vreg_16_10), .down(vreg_16_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_9), .sw(sw));
	wire signed[17:0] vwire_16_10;
	reg signed[17:0] vreg_16_10;
	node n16_10(.left(vreg_15_10), .right(vreg_17_10), .up(vreg_16_11), .down(vreg_16_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_10), .sw(sw));
	wire signed[17:0] vwire_16_11;
	reg signed[17:0] vreg_16_11;
	node n16_11(.left(vreg_15_11), .right(vreg_17_11), .up(vreg_16_12), .down(vreg_16_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_11), .sw(sw));
	wire signed[17:0] vwire_16_12;
	reg signed[17:0] vreg_16_12;
	node n16_12(.left(vreg_15_12), .right(vreg_17_12), .up(vreg_16_13), .down(vreg_16_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_12), .sw(sw));
	wire signed[17:0] vwire_16_13;
	reg signed[17:0] vreg_16_13;
	node n16_13(.left(vreg_15_13), .right(vreg_17_13), .up(vreg_16_14), .down(vreg_16_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_13), .sw(sw));
	wire signed[17:0] vwire_16_14;
	reg signed[17:0] vreg_16_14;
	node n16_14(.left(vreg_15_14), .right(vreg_17_14), .up(vreg_16_15), .down(vreg_16_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_14), .sw(sw));
	wire signed[17:0] vwire_16_15;
	reg signed[17:0] vreg_16_15;
	node n16_15(.left(vreg_15_15), .right(vreg_17_15), .up(vreg_16_16), .down(vreg_16_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_15), .sw(sw));
	wire signed[17:0] vwire_16_16;
	reg signed[17:0] vreg_16_16;
	node n16_16(.left(vreg_15_16), .right(vreg_17_16), .up(vreg_16_17), .down(vreg_16_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_16), .sw(sw));
	wire signed[17:0] vwire_16_17;
	reg signed[17:0] vreg_16_17;
	node n16_17(.left(vreg_15_17), .right(vreg_17_17), .up(vreg_16_18), .down(vreg_16_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_17), .sw(sw));
	wire signed[17:0] vwire_16_18;
	reg signed[17:0] vreg_16_18;
	node n16_18(.left(vreg_15_18), .right(vreg_17_18), .up(vreg_16_19), .down(vreg_16_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_18), .sw(sw));
	wire signed[17:0] vwire_16_19;
	reg signed[17:0] vreg_16_19;
	node n16_19(.left(vreg_15_19), .right(vreg_17_19), .up(vreg_16_20), .down(vreg_16_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_19), .sw(sw));
	wire signed[17:0] vwire_16_20;
	reg signed[17:0] vreg_16_20;
	node n16_20(.left(vreg_15_20), .right(vreg_17_20), .up(vreg_16_21), .down(vreg_16_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_20), .sw(sw));
	wire signed[17:0] vwire_16_21;
	reg signed[17:0] vreg_16_21;
	node n16_21(.left(vreg_15_21), .right(vreg_17_21), .up(vreg_16_22), .down(vreg_16_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_21), .sw(sw));
	wire signed[17:0] vwire_16_22;
	reg signed[17:0] vreg_16_22;
	node n16_22(.left(vreg_15_22), .right(vreg_17_22), .up(vreg_16_23), .down(vreg_16_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_22), .sw(sw));
	wire signed[17:0] vwire_16_23;
	reg signed[17:0] vreg_16_23;
	node n16_23(.left(vreg_15_23), .right(vreg_17_23), .up(vreg_16_24), .down(vreg_16_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_23), .sw(sw));
	wire signed[17:0] vwire_16_24;
	reg signed[17:0] vreg_16_24;
	node n16_24(.left(vreg_15_24), .right(vreg_17_24), .up(vreg_16_25), .down(vreg_16_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_24), .sw(sw));
	wire signed[17:0] vwire_16_25;
	reg signed[17:0] vreg_16_25;
	node n16_25(.left(vreg_15_25), .right(vreg_17_25), .up(vreg_16_26), .down(vreg_16_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_25), .sw(sw));
	wire signed[17:0] vwire_16_26;
	reg signed[17:0] vreg_16_26;
	node n16_26(.left(vreg_15_26), .right(vreg_17_26), .up(vreg_16_27), .down(vreg_16_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_26), .sw(sw));
	wire signed[17:0] vwire_16_27;
	reg signed[17:0] vreg_16_27;
	node n16_27(.left(vreg_15_27), .right(vreg_17_27), .up(vreg_16_28), .down(vreg_16_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_27), .sw(sw));
	wire signed[17:0] vwire_16_28;
	reg signed[17:0] vreg_16_28;
	node n16_28(.left(vreg_15_28), .right(vreg_17_28), .up(vreg_16_29), .down(vreg_16_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_28), .sw(sw));
	wire signed[17:0] vwire_16_29;
	reg signed[17:0] vreg_16_29;
	node n16_29(.left(vreg_15_29), .right(vreg_17_29), .up(vreg_16_30), .down(vreg_16_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_29), .sw(sw));
	wire signed[17:0] vwire_16_30;
	reg signed[17:0] vreg_16_30;
	node n16_30(.left(vreg_15_30), .right(vreg_17_30), .up(vreg_16_31), .down(vreg_16_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_30), .sw(sw));
	wire signed[17:0] vwire_16_31;
	reg signed[17:0] vreg_16_31;
	node n16_31(.left(vreg_15_31), .right(vreg_17_31), .up(vreg_16_32), .down(vreg_16_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_31), .sw(sw));
	wire signed[17:0] vwire_16_32;
	reg signed[17:0] vreg_16_32;
	node n16_32(.left(vreg_15_32), .right(vreg_17_32), .up(vreg_16_33), .down(vreg_16_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_32), .sw(sw));
	wire signed[17:0] vwire_16_33;
	reg signed[17:0] vreg_16_33;
	node n16_33(.left(vreg_15_33), .right(vreg_17_33), .up(vreg_16_34), .down(vreg_16_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_33), .sw(sw));
	wire signed[17:0] vwire_16_34;
	reg signed[17:0] vreg_16_34;
	node n16_34(.left(vreg_15_34), .right(vreg_17_34), .up(vreg_16_35), .down(vreg_16_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_34), .sw(sw));
	wire signed[17:0] vwire_16_35;
	reg signed[17:0] vreg_16_35;
	node n16_35(.left(vreg_15_35), .right(vreg_17_35), .up(vreg_16_36), .down(vreg_16_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_35), .sw(sw));
	wire signed[17:0] vwire_16_36;
	reg signed[17:0] vreg_16_36;
	node n16_36(.left(vreg_15_36), .right(vreg_17_36), .up(vreg_16_37), .down(vreg_16_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_36), .sw(sw));
	wire signed[17:0] vwire_16_37;
	reg signed[17:0] vreg_16_37;
	node n16_37(.left(vreg_15_37), .right(vreg_17_37), .up(vreg_16_38), .down(vreg_16_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_37), .sw(sw));
	wire signed[17:0] vwire_16_38;
	reg signed[17:0] vreg_16_38;
	node n16_38(.left(vreg_15_38), .right(vreg_17_38), .up(vreg_16_39), .down(vreg_16_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_38), .sw(sw));
	wire signed[17:0] vwire_16_39;
	reg signed[17:0] vreg_16_39;
	node n16_39(.left(vreg_15_39), .right(vreg_17_39), .up(vreg_16_40), .down(vreg_16_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_39), .sw(sw));
	wire signed[17:0] vwire_16_40;
	reg signed[17:0] vreg_16_40;
	node n16_40(.left(vreg_15_40), .right(vreg_17_40), .up(vreg_16_41), .down(vreg_16_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_40), .sw(sw));
	wire signed[17:0] vwire_16_41;
	reg signed[17:0] vreg_16_41;
	node n16_41(.left(vreg_15_41), .right(vreg_17_41), .up(vreg_16_42), .down(vreg_16_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_41), .sw(sw));
	wire signed[17:0] vwire_16_42;
	reg signed[17:0] vreg_16_42;
	node n16_42(.left(vreg_15_42), .right(vreg_17_42), .up(vreg_16_43), .down(vreg_16_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_42), .sw(sw));
	wire signed[17:0] vwire_16_43;
	reg signed[17:0] vreg_16_43;
	node n16_43(.left(vreg_15_43), .right(vreg_17_43), .up(vreg_16_44), .down(vreg_16_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_43), .sw(sw));
	wire signed[17:0] vwire_16_44;
	reg signed[17:0] vreg_16_44;
	node n16_44(.left(vreg_15_44), .right(vreg_17_44), .up(vreg_16_45), .down(vreg_16_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_44), .sw(sw));
	wire signed[17:0] vwire_16_45;
	reg signed[17:0] vreg_16_45;
	node n16_45(.left(vreg_15_45), .right(vreg_17_45), .up(vreg_16_46), .down(vreg_16_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_45), .sw(sw));
	wire signed[17:0] vwire_16_46;
	reg signed[17:0] vreg_16_46;
	node n16_46(.left(vreg_15_46), .right(vreg_17_46), .up(vreg_16_47), .down(vreg_16_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_46), .sw(sw));
	wire signed[17:0] vwire_16_47;
	reg signed[17:0] vreg_16_47;
	node n16_47(.left(vreg_15_47), .right(vreg_17_47), .up(vreg_16_48), .down(vreg_16_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_47), .sw(sw));
	wire signed[17:0] vwire_16_48;
	reg signed[17:0] vreg_16_48;
	node n16_48(.left(vreg_15_48), .right(vreg_17_48), .up(vreg_16_49), .down(vreg_16_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_48), .sw(sw));
	wire signed[17:0] vwire_16_49;
	reg signed[17:0] vreg_16_49;
	node n16_49(.left(vreg_15_49), .right(vreg_17_49), .up(18'b0), .down(vreg_16_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_16_49), .sw(sw));
	wire signed[17:0] vwire_17_0;
	reg signed[17:0] vreg_17_0;
	node n17_0(.left(vreg_16_0), .right(vreg_18_0), .up(vreg_17_1), .down(vreg_17_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_0), .sw(sw));
	wire signed[17:0] vwire_17_1;
	reg signed[17:0] vreg_17_1;
	node n17_1(.left(vreg_16_1), .right(vreg_18_1), .up(vreg_17_2), .down(vreg_17_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_1), .sw(sw));
	wire signed[17:0] vwire_17_2;
	reg signed[17:0] vreg_17_2;
	node n17_2(.left(vreg_16_2), .right(vreg_18_2), .up(vreg_17_3), .down(vreg_17_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_2), .sw(sw));
	wire signed[17:0] vwire_17_3;
	reg signed[17:0] vreg_17_3;
	node n17_3(.left(vreg_16_3), .right(vreg_18_3), .up(vreg_17_4), .down(vreg_17_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_3), .sw(sw));
	wire signed[17:0] vwire_17_4;
	reg signed[17:0] vreg_17_4;
	node n17_4(.left(vreg_16_4), .right(vreg_18_4), .up(vreg_17_5), .down(vreg_17_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_4), .sw(sw));
	wire signed[17:0] vwire_17_5;
	reg signed[17:0] vreg_17_5;
	node n17_5(.left(vreg_16_5), .right(vreg_18_5), .up(vreg_17_6), .down(vreg_17_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_5), .sw(sw));
	wire signed[17:0] vwire_17_6;
	reg signed[17:0] vreg_17_6;
	node n17_6(.left(vreg_16_6), .right(vreg_18_6), .up(vreg_17_7), .down(vreg_17_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_6), .sw(sw));
	wire signed[17:0] vwire_17_7;
	reg signed[17:0] vreg_17_7;
	node n17_7(.left(vreg_16_7), .right(vreg_18_7), .up(vreg_17_8), .down(vreg_17_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_7), .sw(sw));
	wire signed[17:0] vwire_17_8;
	reg signed[17:0] vreg_17_8;
	node n17_8(.left(vreg_16_8), .right(vreg_18_8), .up(vreg_17_9), .down(vreg_17_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_8), .sw(sw));
	wire signed[17:0] vwire_17_9;
	reg signed[17:0] vreg_17_9;
	node n17_9(.left(vreg_16_9), .right(vreg_18_9), .up(vreg_17_10), .down(vreg_17_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_9), .sw(sw));
	wire signed[17:0] vwire_17_10;
	reg signed[17:0] vreg_17_10;
	node n17_10(.left(vreg_16_10), .right(vreg_18_10), .up(vreg_17_11), .down(vreg_17_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_10), .sw(sw));
	wire signed[17:0] vwire_17_11;
	reg signed[17:0] vreg_17_11;
	node n17_11(.left(vreg_16_11), .right(vreg_18_11), .up(vreg_17_12), .down(vreg_17_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_11), .sw(sw));
	wire signed[17:0] vwire_17_12;
	reg signed[17:0] vreg_17_12;
	node n17_12(.left(vreg_16_12), .right(vreg_18_12), .up(vreg_17_13), .down(vreg_17_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_12), .sw(sw));
	wire signed[17:0] vwire_17_13;
	reg signed[17:0] vreg_17_13;
	node n17_13(.left(vreg_16_13), .right(vreg_18_13), .up(vreg_17_14), .down(vreg_17_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_13), .sw(sw));
	wire signed[17:0] vwire_17_14;
	reg signed[17:0] vreg_17_14;
	node n17_14(.left(vreg_16_14), .right(vreg_18_14), .up(vreg_17_15), .down(vreg_17_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_14), .sw(sw));
	wire signed[17:0] vwire_17_15;
	reg signed[17:0] vreg_17_15;
	node n17_15(.left(vreg_16_15), .right(vreg_18_15), .up(vreg_17_16), .down(vreg_17_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_15), .sw(sw));
	wire signed[17:0] vwire_17_16;
	reg signed[17:0] vreg_17_16;
	node n17_16(.left(vreg_16_16), .right(vreg_18_16), .up(vreg_17_17), .down(vreg_17_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_16), .sw(sw));
	wire signed[17:0] vwire_17_17;
	reg signed[17:0] vreg_17_17;
	node n17_17(.left(vreg_16_17), .right(vreg_18_17), .up(vreg_17_18), .down(vreg_17_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_17), .sw(sw));
	wire signed[17:0] vwire_17_18;
	reg signed[17:0] vreg_17_18;
	node n17_18(.left(vreg_16_18), .right(vreg_18_18), .up(vreg_17_19), .down(vreg_17_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_18), .sw(sw));
	wire signed[17:0] vwire_17_19;
	reg signed[17:0] vreg_17_19;
	node n17_19(.left(vreg_16_19), .right(vreg_18_19), .up(vreg_17_20), .down(vreg_17_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_19), .sw(sw));
	wire signed[17:0] vwire_17_20;
	reg signed[17:0] vreg_17_20;
	node n17_20(.left(vreg_16_20), .right(vreg_18_20), .up(vreg_17_21), .down(vreg_17_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_20), .sw(sw));
	wire signed[17:0] vwire_17_21;
	reg signed[17:0] vreg_17_21;
	node n17_21(.left(vreg_16_21), .right(vreg_18_21), .up(vreg_17_22), .down(vreg_17_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_21), .sw(sw));
	wire signed[17:0] vwire_17_22;
	reg signed[17:0] vreg_17_22;
	node n17_22(.left(vreg_16_22), .right(vreg_18_22), .up(vreg_17_23), .down(vreg_17_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_22), .sw(sw));
	wire signed[17:0] vwire_17_23;
	reg signed[17:0] vreg_17_23;
	node n17_23(.left(vreg_16_23), .right(vreg_18_23), .up(vreg_17_24), .down(vreg_17_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_23), .sw(sw));
	wire signed[17:0] vwire_17_24;
	reg signed[17:0] vreg_17_24;
	node n17_24(.left(vreg_16_24), .right(vreg_18_24), .up(vreg_17_25), .down(vreg_17_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_24), .sw(sw));
	wire signed[17:0] vwire_17_25;
	reg signed[17:0] vreg_17_25;
	node n17_25(.left(vreg_16_25), .right(vreg_18_25), .up(vreg_17_26), .down(vreg_17_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_25), .sw(sw));
	wire signed[17:0] vwire_17_26;
	reg signed[17:0] vreg_17_26;
	node n17_26(.left(vreg_16_26), .right(vreg_18_26), .up(vreg_17_27), .down(vreg_17_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_26), .sw(sw));
	wire signed[17:0] vwire_17_27;
	reg signed[17:0] vreg_17_27;
	node n17_27(.left(vreg_16_27), .right(vreg_18_27), .up(vreg_17_28), .down(vreg_17_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_27), .sw(sw));
	wire signed[17:0] vwire_17_28;
	reg signed[17:0] vreg_17_28;
	node n17_28(.left(vreg_16_28), .right(vreg_18_28), .up(vreg_17_29), .down(vreg_17_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_28), .sw(sw));
	wire signed[17:0] vwire_17_29;
	reg signed[17:0] vreg_17_29;
	node n17_29(.left(vreg_16_29), .right(vreg_18_29), .up(vreg_17_30), .down(vreg_17_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_29), .sw(sw));
	wire signed[17:0] vwire_17_30;
	reg signed[17:0] vreg_17_30;
	node n17_30(.left(vreg_16_30), .right(vreg_18_30), .up(vreg_17_31), .down(vreg_17_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_30), .sw(sw));
	wire signed[17:0] vwire_17_31;
	reg signed[17:0] vreg_17_31;
	node n17_31(.left(vreg_16_31), .right(vreg_18_31), .up(vreg_17_32), .down(vreg_17_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_31), .sw(sw));
	wire signed[17:0] vwire_17_32;
	reg signed[17:0] vreg_17_32;
	node n17_32(.left(vreg_16_32), .right(vreg_18_32), .up(vreg_17_33), .down(vreg_17_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_32), .sw(sw));
	wire signed[17:0] vwire_17_33;
	reg signed[17:0] vreg_17_33;
	node n17_33(.left(vreg_16_33), .right(vreg_18_33), .up(vreg_17_34), .down(vreg_17_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_33), .sw(sw));
	wire signed[17:0] vwire_17_34;
	reg signed[17:0] vreg_17_34;
	node n17_34(.left(vreg_16_34), .right(vreg_18_34), .up(vreg_17_35), .down(vreg_17_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_34), .sw(sw));
	wire signed[17:0] vwire_17_35;
	reg signed[17:0] vreg_17_35;
	node n17_35(.left(vreg_16_35), .right(vreg_18_35), .up(vreg_17_36), .down(vreg_17_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_35), .sw(sw));
	wire signed[17:0] vwire_17_36;
	reg signed[17:0] vreg_17_36;
	node n17_36(.left(vreg_16_36), .right(vreg_18_36), .up(vreg_17_37), .down(vreg_17_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_36), .sw(sw));
	wire signed[17:0] vwire_17_37;
	reg signed[17:0] vreg_17_37;
	node n17_37(.left(vreg_16_37), .right(vreg_18_37), .up(vreg_17_38), .down(vreg_17_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_37), .sw(sw));
	wire signed[17:0] vwire_17_38;
	reg signed[17:0] vreg_17_38;
	node n17_38(.left(vreg_16_38), .right(vreg_18_38), .up(vreg_17_39), .down(vreg_17_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_38), .sw(sw));
	wire signed[17:0] vwire_17_39;
	reg signed[17:0] vreg_17_39;
	node n17_39(.left(vreg_16_39), .right(vreg_18_39), .up(vreg_17_40), .down(vreg_17_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_39), .sw(sw));
	wire signed[17:0] vwire_17_40;
	reg signed[17:0] vreg_17_40;
	node n17_40(.left(vreg_16_40), .right(vreg_18_40), .up(vreg_17_41), .down(vreg_17_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_40), .sw(sw));
	wire signed[17:0] vwire_17_41;
	reg signed[17:0] vreg_17_41;
	node n17_41(.left(vreg_16_41), .right(vreg_18_41), .up(vreg_17_42), .down(vreg_17_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_41), .sw(sw));
	wire signed[17:0] vwire_17_42;
	reg signed[17:0] vreg_17_42;
	node n17_42(.left(vreg_16_42), .right(vreg_18_42), .up(vreg_17_43), .down(vreg_17_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_42), .sw(sw));
	wire signed[17:0] vwire_17_43;
	reg signed[17:0] vreg_17_43;
	node n17_43(.left(vreg_16_43), .right(vreg_18_43), .up(vreg_17_44), .down(vreg_17_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_43), .sw(sw));
	wire signed[17:0] vwire_17_44;
	reg signed[17:0] vreg_17_44;
	node n17_44(.left(vreg_16_44), .right(vreg_18_44), .up(vreg_17_45), .down(vreg_17_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_44), .sw(sw));
	wire signed[17:0] vwire_17_45;
	reg signed[17:0] vreg_17_45;
	node n17_45(.left(vreg_16_45), .right(vreg_18_45), .up(vreg_17_46), .down(vreg_17_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_45), .sw(sw));
	wire signed[17:0] vwire_17_46;
	reg signed[17:0] vreg_17_46;
	node n17_46(.left(vreg_16_46), .right(vreg_18_46), .up(vreg_17_47), .down(vreg_17_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_46), .sw(sw));
	wire signed[17:0] vwire_17_47;
	reg signed[17:0] vreg_17_47;
	node n17_47(.left(vreg_16_47), .right(vreg_18_47), .up(vreg_17_48), .down(vreg_17_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_47), .sw(sw));
	wire signed[17:0] vwire_17_48;
	reg signed[17:0] vreg_17_48;
	node n17_48(.left(vreg_16_48), .right(vreg_18_48), .up(vreg_17_49), .down(vreg_17_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_48), .sw(sw));
	wire signed[17:0] vwire_17_49;
	reg signed[17:0] vreg_17_49;
	node n17_49(.left(vreg_16_49), .right(vreg_18_49), .up(18'b0), .down(vreg_17_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_17_49), .sw(sw));
	wire signed[17:0] vwire_18_0;
	reg signed[17:0] vreg_18_0;
	node n18_0(.left(vreg_17_0), .right(vreg_19_0), .up(vreg_18_1), .down(vreg_18_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_0), .sw(sw));
	wire signed[17:0] vwire_18_1;
	reg signed[17:0] vreg_18_1;
	node n18_1(.left(vreg_17_1), .right(vreg_19_1), .up(vreg_18_2), .down(vreg_18_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_1), .sw(sw));
	wire signed[17:0] vwire_18_2;
	reg signed[17:0] vreg_18_2;
	node n18_2(.left(vreg_17_2), .right(vreg_19_2), .up(vreg_18_3), .down(vreg_18_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_2), .sw(sw));
	wire signed[17:0] vwire_18_3;
	reg signed[17:0] vreg_18_3;
	node n18_3(.left(vreg_17_3), .right(vreg_19_3), .up(vreg_18_4), .down(vreg_18_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_3), .sw(sw));
	wire signed[17:0] vwire_18_4;
	reg signed[17:0] vreg_18_4;
	node n18_4(.left(vreg_17_4), .right(vreg_19_4), .up(vreg_18_5), .down(vreg_18_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_4), .sw(sw));
	wire signed[17:0] vwire_18_5;
	reg signed[17:0] vreg_18_5;
	node n18_5(.left(vreg_17_5), .right(vreg_19_5), .up(vreg_18_6), .down(vreg_18_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_5), .sw(sw));
	wire signed[17:0] vwire_18_6;
	reg signed[17:0] vreg_18_6;
	node n18_6(.left(vreg_17_6), .right(vreg_19_6), .up(vreg_18_7), .down(vreg_18_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_6), .sw(sw));
	wire signed[17:0] vwire_18_7;
	reg signed[17:0] vreg_18_7;
	node n18_7(.left(vreg_17_7), .right(vreg_19_7), .up(vreg_18_8), .down(vreg_18_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_7), .sw(sw));
	wire signed[17:0] vwire_18_8;
	reg signed[17:0] vreg_18_8;
	node n18_8(.left(vreg_17_8), .right(vreg_19_8), .up(vreg_18_9), .down(vreg_18_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_8), .sw(sw));
	wire signed[17:0] vwire_18_9;
	reg signed[17:0] vreg_18_9;
	node n18_9(.left(vreg_17_9), .right(vreg_19_9), .up(vreg_18_10), .down(vreg_18_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_9), .sw(sw));
	wire signed[17:0] vwire_18_10;
	reg signed[17:0] vreg_18_10;
	node n18_10(.left(vreg_17_10), .right(vreg_19_10), .up(vreg_18_11), .down(vreg_18_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_10), .sw(sw));
	wire signed[17:0] vwire_18_11;
	reg signed[17:0] vreg_18_11;
	node n18_11(.left(vreg_17_11), .right(vreg_19_11), .up(vreg_18_12), .down(vreg_18_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_11), .sw(sw));
	wire signed[17:0] vwire_18_12;
	reg signed[17:0] vreg_18_12;
	node n18_12(.left(vreg_17_12), .right(vreg_19_12), .up(vreg_18_13), .down(vreg_18_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_12), .sw(sw));
	wire signed[17:0] vwire_18_13;
	reg signed[17:0] vreg_18_13;
	node n18_13(.left(vreg_17_13), .right(vreg_19_13), .up(vreg_18_14), .down(vreg_18_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_13), .sw(sw));
	wire signed[17:0] vwire_18_14;
	reg signed[17:0] vreg_18_14;
	node n18_14(.left(vreg_17_14), .right(vreg_19_14), .up(vreg_18_15), .down(vreg_18_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_14), .sw(sw));
	wire signed[17:0] vwire_18_15;
	reg signed[17:0] vreg_18_15;
	node n18_15(.left(vreg_17_15), .right(vreg_19_15), .up(vreg_18_16), .down(vreg_18_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_15), .sw(sw));
	wire signed[17:0] vwire_18_16;
	reg signed[17:0] vreg_18_16;
	node n18_16(.left(vreg_17_16), .right(vreg_19_16), .up(vreg_18_17), .down(vreg_18_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_16), .sw(sw));
	wire signed[17:0] vwire_18_17;
	reg signed[17:0] vreg_18_17;
	node n18_17(.left(vreg_17_17), .right(vreg_19_17), .up(vreg_18_18), .down(vreg_18_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_17), .sw(sw));
	wire signed[17:0] vwire_18_18;
	reg signed[17:0] vreg_18_18;
	node n18_18(.left(vreg_17_18), .right(vreg_19_18), .up(vreg_18_19), .down(vreg_18_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_18), .sw(sw));
	wire signed[17:0] vwire_18_19;
	reg signed[17:0] vreg_18_19;
	node n18_19(.left(vreg_17_19), .right(vreg_19_19), .up(vreg_18_20), .down(vreg_18_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_19), .sw(sw));
	wire signed[17:0] vwire_18_20;
	reg signed[17:0] vreg_18_20;
	node n18_20(.left(vreg_17_20), .right(vreg_19_20), .up(vreg_18_21), .down(vreg_18_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_20), .sw(sw));
	wire signed[17:0] vwire_18_21;
	reg signed[17:0] vreg_18_21;
	node n18_21(.left(vreg_17_21), .right(vreg_19_21), .up(vreg_18_22), .down(vreg_18_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_21), .sw(sw));
	wire signed[17:0] vwire_18_22;
	reg signed[17:0] vreg_18_22;
	node n18_22(.left(vreg_17_22), .right(vreg_19_22), .up(vreg_18_23), .down(vreg_18_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_22), .sw(sw));
	wire signed[17:0] vwire_18_23;
	reg signed[17:0] vreg_18_23;
	node n18_23(.left(vreg_17_23), .right(vreg_19_23), .up(vreg_18_24), .down(vreg_18_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_23), .sw(sw));
	wire signed[17:0] vwire_18_24;
	reg signed[17:0] vreg_18_24;
	node n18_24(.left(vreg_17_24), .right(vreg_19_24), .up(vreg_18_25), .down(vreg_18_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_24), .sw(sw));
	wire signed[17:0] vwire_18_25;
	reg signed[17:0] vreg_18_25;
	node n18_25(.left(vreg_17_25), .right(vreg_19_25), .up(vreg_18_26), .down(vreg_18_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_25), .sw(sw));
	wire signed[17:0] vwire_18_26;
	reg signed[17:0] vreg_18_26;
	node n18_26(.left(vreg_17_26), .right(vreg_19_26), .up(vreg_18_27), .down(vreg_18_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_26), .sw(sw));
	wire signed[17:0] vwire_18_27;
	reg signed[17:0] vreg_18_27;
	node n18_27(.left(vreg_17_27), .right(vreg_19_27), .up(vreg_18_28), .down(vreg_18_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_27), .sw(sw));
	wire signed[17:0] vwire_18_28;
	reg signed[17:0] vreg_18_28;
	node n18_28(.left(vreg_17_28), .right(vreg_19_28), .up(vreg_18_29), .down(vreg_18_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_28), .sw(sw));
	wire signed[17:0] vwire_18_29;
	reg signed[17:0] vreg_18_29;
	node n18_29(.left(vreg_17_29), .right(vreg_19_29), .up(vreg_18_30), .down(vreg_18_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_29), .sw(sw));
	wire signed[17:0] vwire_18_30;
	reg signed[17:0] vreg_18_30;
	node n18_30(.left(vreg_17_30), .right(vreg_19_30), .up(vreg_18_31), .down(vreg_18_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_30), .sw(sw));
	wire signed[17:0] vwire_18_31;
	reg signed[17:0] vreg_18_31;
	node n18_31(.left(vreg_17_31), .right(vreg_19_31), .up(vreg_18_32), .down(vreg_18_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_31), .sw(sw));
	wire signed[17:0] vwire_18_32;
	reg signed[17:0] vreg_18_32;
	node n18_32(.left(vreg_17_32), .right(vreg_19_32), .up(vreg_18_33), .down(vreg_18_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_32), .sw(sw));
	wire signed[17:0] vwire_18_33;
	reg signed[17:0] vreg_18_33;
	node n18_33(.left(vreg_17_33), .right(vreg_19_33), .up(vreg_18_34), .down(vreg_18_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_33), .sw(sw));
	wire signed[17:0] vwire_18_34;
	reg signed[17:0] vreg_18_34;
	node n18_34(.left(vreg_17_34), .right(vreg_19_34), .up(vreg_18_35), .down(vreg_18_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_34), .sw(sw));
	wire signed[17:0] vwire_18_35;
	reg signed[17:0] vreg_18_35;
	node n18_35(.left(vreg_17_35), .right(vreg_19_35), .up(vreg_18_36), .down(vreg_18_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_35), .sw(sw));
	wire signed[17:0] vwire_18_36;
	reg signed[17:0] vreg_18_36;
	node n18_36(.left(vreg_17_36), .right(vreg_19_36), .up(vreg_18_37), .down(vreg_18_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_36), .sw(sw));
	wire signed[17:0] vwire_18_37;
	reg signed[17:0] vreg_18_37;
	node n18_37(.left(vreg_17_37), .right(vreg_19_37), .up(vreg_18_38), .down(vreg_18_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_37), .sw(sw));
	wire signed[17:0] vwire_18_38;
	reg signed[17:0] vreg_18_38;
	node n18_38(.left(vreg_17_38), .right(vreg_19_38), .up(vreg_18_39), .down(vreg_18_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_38), .sw(sw));
	wire signed[17:0] vwire_18_39;
	reg signed[17:0] vreg_18_39;
	node n18_39(.left(vreg_17_39), .right(vreg_19_39), .up(vreg_18_40), .down(vreg_18_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_39), .sw(sw));
	wire signed[17:0] vwire_18_40;
	reg signed[17:0] vreg_18_40;
	node n18_40(.left(vreg_17_40), .right(vreg_19_40), .up(vreg_18_41), .down(vreg_18_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_40), .sw(sw));
	wire signed[17:0] vwire_18_41;
	reg signed[17:0] vreg_18_41;
	node n18_41(.left(vreg_17_41), .right(vreg_19_41), .up(vreg_18_42), .down(vreg_18_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_41), .sw(sw));
	wire signed[17:0] vwire_18_42;
	reg signed[17:0] vreg_18_42;
	node n18_42(.left(vreg_17_42), .right(vreg_19_42), .up(vreg_18_43), .down(vreg_18_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_42), .sw(sw));
	wire signed[17:0] vwire_18_43;
	reg signed[17:0] vreg_18_43;
	node n18_43(.left(vreg_17_43), .right(vreg_19_43), .up(vreg_18_44), .down(vreg_18_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_43), .sw(sw));
	wire signed[17:0] vwire_18_44;
	reg signed[17:0] vreg_18_44;
	node n18_44(.left(vreg_17_44), .right(vreg_19_44), .up(vreg_18_45), .down(vreg_18_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_44), .sw(sw));
	wire signed[17:0] vwire_18_45;
	reg signed[17:0] vreg_18_45;
	node n18_45(.left(vreg_17_45), .right(vreg_19_45), .up(vreg_18_46), .down(vreg_18_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_45), .sw(sw));
	wire signed[17:0] vwire_18_46;
	reg signed[17:0] vreg_18_46;
	node n18_46(.left(vreg_17_46), .right(vreg_19_46), .up(vreg_18_47), .down(vreg_18_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_46), .sw(sw));
	wire signed[17:0] vwire_18_47;
	reg signed[17:0] vreg_18_47;
	node n18_47(.left(vreg_17_47), .right(vreg_19_47), .up(vreg_18_48), .down(vreg_18_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_47), .sw(sw));
	wire signed[17:0] vwire_18_48;
	reg signed[17:0] vreg_18_48;
	node n18_48(.left(vreg_17_48), .right(vreg_19_48), .up(vreg_18_49), .down(vreg_18_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_48), .sw(sw));
	wire signed[17:0] vwire_18_49;
	reg signed[17:0] vreg_18_49;
	node n18_49(.left(vreg_17_49), .right(vreg_19_49), .up(18'b0), .down(vreg_18_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_18_49), .sw(sw));
	wire signed[17:0] vwire_19_0;
	reg signed[17:0] vreg_19_0;
	node n19_0(.left(vreg_18_0), .right(vreg_20_0), .up(vreg_19_1), .down(vreg_19_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_0), .sw(sw));
	wire signed[17:0] vwire_19_1;
	reg signed[17:0] vreg_19_1;
	node n19_1(.left(vreg_18_1), .right(vreg_20_1), .up(vreg_19_2), .down(vreg_19_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_1), .sw(sw));
	wire signed[17:0] vwire_19_2;
	reg signed[17:0] vreg_19_2;
	node n19_2(.left(vreg_18_2), .right(vreg_20_2), .up(vreg_19_3), .down(vreg_19_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_2), .sw(sw));
	wire signed[17:0] vwire_19_3;
	reg signed[17:0] vreg_19_3;
	node n19_3(.left(vreg_18_3), .right(vreg_20_3), .up(vreg_19_4), .down(vreg_19_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_3), .sw(sw));
	wire signed[17:0] vwire_19_4;
	reg signed[17:0] vreg_19_4;
	node n19_4(.left(vreg_18_4), .right(vreg_20_4), .up(vreg_19_5), .down(vreg_19_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_4), .sw(sw));
	wire signed[17:0] vwire_19_5;
	reg signed[17:0] vreg_19_5;
	node n19_5(.left(vreg_18_5), .right(vreg_20_5), .up(vreg_19_6), .down(vreg_19_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_5), .sw(sw));
	wire signed[17:0] vwire_19_6;
	reg signed[17:0] vreg_19_6;
	node n19_6(.left(vreg_18_6), .right(vreg_20_6), .up(vreg_19_7), .down(vreg_19_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_6), .sw(sw));
	wire signed[17:0] vwire_19_7;
	reg signed[17:0] vreg_19_7;
	node n19_7(.left(vreg_18_7), .right(vreg_20_7), .up(vreg_19_8), .down(vreg_19_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_7), .sw(sw));
	wire signed[17:0] vwire_19_8;
	reg signed[17:0] vreg_19_8;
	node n19_8(.left(vreg_18_8), .right(vreg_20_8), .up(vreg_19_9), .down(vreg_19_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_8), .sw(sw));
	wire signed[17:0] vwire_19_9;
	reg signed[17:0] vreg_19_9;
	node n19_9(.left(vreg_18_9), .right(vreg_20_9), .up(vreg_19_10), .down(vreg_19_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_9), .sw(sw));
	wire signed[17:0] vwire_19_10;
	reg signed[17:0] vreg_19_10;
	node n19_10(.left(vreg_18_10), .right(vreg_20_10), .up(vreg_19_11), .down(vreg_19_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_10), .sw(sw));
	wire signed[17:0] vwire_19_11;
	reg signed[17:0] vreg_19_11;
	node n19_11(.left(vreg_18_11), .right(vreg_20_11), .up(vreg_19_12), .down(vreg_19_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_11), .sw(sw));
	wire signed[17:0] vwire_19_12;
	reg signed[17:0] vreg_19_12;
	node n19_12(.left(vreg_18_12), .right(vreg_20_12), .up(vreg_19_13), .down(vreg_19_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_12), .sw(sw));
	wire signed[17:0] vwire_19_13;
	reg signed[17:0] vreg_19_13;
	node n19_13(.left(vreg_18_13), .right(vreg_20_13), .up(vreg_19_14), .down(vreg_19_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_13), .sw(sw));
	wire signed[17:0] vwire_19_14;
	reg signed[17:0] vreg_19_14;
	node n19_14(.left(vreg_18_14), .right(vreg_20_14), .up(vreg_19_15), .down(vreg_19_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_14), .sw(sw));
	wire signed[17:0] vwire_19_15;
	reg signed[17:0] vreg_19_15;
	node n19_15(.left(vreg_18_15), .right(vreg_20_15), .up(vreg_19_16), .down(vreg_19_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_15), .sw(sw));
	wire signed[17:0] vwire_19_16;
	reg signed[17:0] vreg_19_16;
	node n19_16(.left(vreg_18_16), .right(vreg_20_16), .up(vreg_19_17), .down(vreg_19_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_16), .sw(sw));
	wire signed[17:0] vwire_19_17;
	reg signed[17:0] vreg_19_17;
	node n19_17(.left(vreg_18_17), .right(vreg_20_17), .up(vreg_19_18), .down(vreg_19_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_17), .sw(sw));
	wire signed[17:0] vwire_19_18;
	reg signed[17:0] vreg_19_18;
	node n19_18(.left(vreg_18_18), .right(vreg_20_18), .up(vreg_19_19), .down(vreg_19_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_18), .sw(sw));
	wire signed[17:0] vwire_19_19;
	reg signed[17:0] vreg_19_19;
	node n19_19(.left(vreg_18_19), .right(vreg_20_19), .up(vreg_19_20), .down(vreg_19_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_19), .sw(sw));
	wire signed[17:0] vwire_19_20;
	reg signed[17:0] vreg_19_20;
	node n19_20(.left(vreg_18_20), .right(vreg_20_20), .up(vreg_19_21), .down(vreg_19_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_20), .sw(sw));
	wire signed[17:0] vwire_19_21;
	reg signed[17:0] vreg_19_21;
	node n19_21(.left(vreg_18_21), .right(vreg_20_21), .up(vreg_19_22), .down(vreg_19_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_21), .sw(sw));
	wire signed[17:0] vwire_19_22;
	reg signed[17:0] vreg_19_22;
	node n19_22(.left(vreg_18_22), .right(vreg_20_22), .up(vreg_19_23), .down(vreg_19_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_22), .sw(sw));
	wire signed[17:0] vwire_19_23;
	reg signed[17:0] vreg_19_23;
	node n19_23(.left(vreg_18_23), .right(vreg_20_23), .up(vreg_19_24), .down(vreg_19_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_23), .sw(sw));
	wire signed[17:0] vwire_19_24;
	reg signed[17:0] vreg_19_24;
	node n19_24(.left(vreg_18_24), .right(vreg_20_24), .up(vreg_19_25), .down(vreg_19_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_24), .sw(sw));
	wire signed[17:0] vwire_19_25;
	reg signed[17:0] vreg_19_25;
	node n19_25(.left(vreg_18_25), .right(vreg_20_25), .up(vreg_19_26), .down(vreg_19_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_25), .sw(sw));
	wire signed[17:0] vwire_19_26;
	reg signed[17:0] vreg_19_26;
	node n19_26(.left(vreg_18_26), .right(vreg_20_26), .up(vreg_19_27), .down(vreg_19_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_26), .sw(sw));
	wire signed[17:0] vwire_19_27;
	reg signed[17:0] vreg_19_27;
	node n19_27(.left(vreg_18_27), .right(vreg_20_27), .up(vreg_19_28), .down(vreg_19_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_27), .sw(sw));
	wire signed[17:0] vwire_19_28;
	reg signed[17:0] vreg_19_28;
	node n19_28(.left(vreg_18_28), .right(vreg_20_28), .up(vreg_19_29), .down(vreg_19_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_28), .sw(sw));
	wire signed[17:0] vwire_19_29;
	reg signed[17:0] vreg_19_29;
	node n19_29(.left(vreg_18_29), .right(vreg_20_29), .up(vreg_19_30), .down(vreg_19_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_29), .sw(sw));
	wire signed[17:0] vwire_19_30;
	reg signed[17:0] vreg_19_30;
	node n19_30(.left(vreg_18_30), .right(vreg_20_30), .up(vreg_19_31), .down(vreg_19_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_30), .sw(sw));
	wire signed[17:0] vwire_19_31;
	reg signed[17:0] vreg_19_31;
	node n19_31(.left(vreg_18_31), .right(vreg_20_31), .up(vreg_19_32), .down(vreg_19_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_31), .sw(sw));
	wire signed[17:0] vwire_19_32;
	reg signed[17:0] vreg_19_32;
	node n19_32(.left(vreg_18_32), .right(vreg_20_32), .up(vreg_19_33), .down(vreg_19_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_32), .sw(sw));
	wire signed[17:0] vwire_19_33;
	reg signed[17:0] vreg_19_33;
	node n19_33(.left(vreg_18_33), .right(vreg_20_33), .up(vreg_19_34), .down(vreg_19_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_33), .sw(sw));
	wire signed[17:0] vwire_19_34;
	reg signed[17:0] vreg_19_34;
	node n19_34(.left(vreg_18_34), .right(vreg_20_34), .up(vreg_19_35), .down(vreg_19_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_34), .sw(sw));
	wire signed[17:0] vwire_19_35;
	reg signed[17:0] vreg_19_35;
	node n19_35(.left(vreg_18_35), .right(vreg_20_35), .up(vreg_19_36), .down(vreg_19_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_35), .sw(sw));
	wire signed[17:0] vwire_19_36;
	reg signed[17:0] vreg_19_36;
	node n19_36(.left(vreg_18_36), .right(vreg_20_36), .up(vreg_19_37), .down(vreg_19_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_36), .sw(sw));
	wire signed[17:0] vwire_19_37;
	reg signed[17:0] vreg_19_37;
	node n19_37(.left(vreg_18_37), .right(vreg_20_37), .up(vreg_19_38), .down(vreg_19_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_37), .sw(sw));
	wire signed[17:0] vwire_19_38;
	reg signed[17:0] vreg_19_38;
	node n19_38(.left(vreg_18_38), .right(vreg_20_38), .up(vreg_19_39), .down(vreg_19_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_38), .sw(sw));
	wire signed[17:0] vwire_19_39;
	reg signed[17:0] vreg_19_39;
	node n19_39(.left(vreg_18_39), .right(vreg_20_39), .up(vreg_19_40), .down(vreg_19_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_39), .sw(sw));
	wire signed[17:0] vwire_19_40;
	reg signed[17:0] vreg_19_40;
	node n19_40(.left(vreg_18_40), .right(vreg_20_40), .up(vreg_19_41), .down(vreg_19_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_40), .sw(sw));
	wire signed[17:0] vwire_19_41;
	reg signed[17:0] vreg_19_41;
	node n19_41(.left(vreg_18_41), .right(vreg_20_41), .up(vreg_19_42), .down(vreg_19_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_41), .sw(sw));
	wire signed[17:0] vwire_19_42;
	reg signed[17:0] vreg_19_42;
	node n19_42(.left(vreg_18_42), .right(vreg_20_42), .up(vreg_19_43), .down(vreg_19_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_42), .sw(sw));
	wire signed[17:0] vwire_19_43;
	reg signed[17:0] vreg_19_43;
	node n19_43(.left(vreg_18_43), .right(vreg_20_43), .up(vreg_19_44), .down(vreg_19_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_43), .sw(sw));
	wire signed[17:0] vwire_19_44;
	reg signed[17:0] vreg_19_44;
	node n19_44(.left(vreg_18_44), .right(vreg_20_44), .up(vreg_19_45), .down(vreg_19_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_44), .sw(sw));
	wire signed[17:0] vwire_19_45;
	reg signed[17:0] vreg_19_45;
	node n19_45(.left(vreg_18_45), .right(vreg_20_45), .up(vreg_19_46), .down(vreg_19_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_45), .sw(sw));
	wire signed[17:0] vwire_19_46;
	reg signed[17:0] vreg_19_46;
	node n19_46(.left(vreg_18_46), .right(vreg_20_46), .up(vreg_19_47), .down(vreg_19_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_46), .sw(sw));
	wire signed[17:0] vwire_19_47;
	reg signed[17:0] vreg_19_47;
	node n19_47(.left(vreg_18_47), .right(vreg_20_47), .up(vreg_19_48), .down(vreg_19_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_47), .sw(sw));
	wire signed[17:0] vwire_19_48;
	reg signed[17:0] vreg_19_48;
	node n19_48(.left(vreg_18_48), .right(vreg_20_48), .up(vreg_19_49), .down(vreg_19_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_48), .sw(sw));
	wire signed[17:0] vwire_19_49;
	reg signed[17:0] vreg_19_49;
	node n19_49(.left(vreg_18_49), .right(vreg_20_49), .up(18'b0), .down(vreg_19_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_19_49), .sw(sw));
	wire signed[17:0] vwire_20_0;
	reg signed[17:0] vreg_20_0;
	node n20_0(.left(vreg_19_0), .right(vreg_21_0), .up(vreg_20_1), .down(vreg_20_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_0), .sw(sw));
	wire signed[17:0] vwire_20_1;
	reg signed[17:0] vreg_20_1;
	node n20_1(.left(vreg_19_1), .right(vreg_21_1), .up(vreg_20_2), .down(vreg_20_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_1), .sw(sw));
	wire signed[17:0] vwire_20_2;
	reg signed[17:0] vreg_20_2;
	node n20_2(.left(vreg_19_2), .right(vreg_21_2), .up(vreg_20_3), .down(vreg_20_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_2), .sw(sw));
	wire signed[17:0] vwire_20_3;
	reg signed[17:0] vreg_20_3;
	node n20_3(.left(vreg_19_3), .right(vreg_21_3), .up(vreg_20_4), .down(vreg_20_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_3), .sw(sw));
	wire signed[17:0] vwire_20_4;
	reg signed[17:0] vreg_20_4;
	node n20_4(.left(vreg_19_4), .right(vreg_21_4), .up(vreg_20_5), .down(vreg_20_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_4), .sw(sw));
	wire signed[17:0] vwire_20_5;
	reg signed[17:0] vreg_20_5;
	node n20_5(.left(vreg_19_5), .right(vreg_21_5), .up(vreg_20_6), .down(vreg_20_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_5), .sw(sw));
	wire signed[17:0] vwire_20_6;
	reg signed[17:0] vreg_20_6;
	node n20_6(.left(vreg_19_6), .right(vreg_21_6), .up(vreg_20_7), .down(vreg_20_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_6), .sw(sw));
	wire signed[17:0] vwire_20_7;
	reg signed[17:0] vreg_20_7;
	node n20_7(.left(vreg_19_7), .right(vreg_21_7), .up(vreg_20_8), .down(vreg_20_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_7), .sw(sw));
	wire signed[17:0] vwire_20_8;
	reg signed[17:0] vreg_20_8;
	node n20_8(.left(vreg_19_8), .right(vreg_21_8), .up(vreg_20_9), .down(vreg_20_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_8), .sw(sw));
	wire signed[17:0] vwire_20_9;
	reg signed[17:0] vreg_20_9;
	node n20_9(.left(vreg_19_9), .right(vreg_21_9), .up(vreg_20_10), .down(vreg_20_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_9), .sw(sw));
	wire signed[17:0] vwire_20_10;
	reg signed[17:0] vreg_20_10;
	node n20_10(.left(vreg_19_10), .right(vreg_21_10), .up(vreg_20_11), .down(vreg_20_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_10), .sw(sw));
	wire signed[17:0] vwire_20_11;
	reg signed[17:0] vreg_20_11;
	node n20_11(.left(vreg_19_11), .right(vreg_21_11), .up(vreg_20_12), .down(vreg_20_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_11), .sw(sw));
	wire signed[17:0] vwire_20_12;
	reg signed[17:0] vreg_20_12;
	node n20_12(.left(vreg_19_12), .right(vreg_21_12), .up(vreg_20_13), .down(vreg_20_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_12), .sw(sw));
	wire signed[17:0] vwire_20_13;
	reg signed[17:0] vreg_20_13;
	node n20_13(.left(vreg_19_13), .right(vreg_21_13), .up(vreg_20_14), .down(vreg_20_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_13), .sw(sw));
	wire signed[17:0] vwire_20_14;
	reg signed[17:0] vreg_20_14;
	node n20_14(.left(vreg_19_14), .right(vreg_21_14), .up(vreg_20_15), .down(vreg_20_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_14), .sw(sw));
	wire signed[17:0] vwire_20_15;
	reg signed[17:0] vreg_20_15;
	node n20_15(.left(vreg_19_15), .right(vreg_21_15), .up(vreg_20_16), .down(vreg_20_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_15), .sw(sw));
	wire signed[17:0] vwire_20_16;
	reg signed[17:0] vreg_20_16;
	node n20_16(.left(vreg_19_16), .right(vreg_21_16), .up(vreg_20_17), .down(vreg_20_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_16), .sw(sw));
	wire signed[17:0] vwire_20_17;
	reg signed[17:0] vreg_20_17;
	node n20_17(.left(vreg_19_17), .right(vreg_21_17), .up(vreg_20_18), .down(vreg_20_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_17), .sw(sw));
	wire signed[17:0] vwire_20_18;
	reg signed[17:0] vreg_20_18;
	node n20_18(.left(vreg_19_18), .right(vreg_21_18), .up(vreg_20_19), .down(vreg_20_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_18), .sw(sw));
	wire signed[17:0] vwire_20_19;
	reg signed[17:0] vreg_20_19;
	node n20_19(.left(vreg_19_19), .right(vreg_21_19), .up(vreg_20_20), .down(vreg_20_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_19), .sw(sw));
	wire signed[17:0] vwire_20_20;
	reg signed[17:0] vreg_20_20;
	node n20_20(.left(vreg_19_20), .right(vreg_21_20), .up(vreg_20_21), .down(vreg_20_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_20), .sw(sw));
	wire signed[17:0] vwire_20_21;
	reg signed[17:0] vreg_20_21;
	node n20_21(.left(vreg_19_21), .right(vreg_21_21), .up(vreg_20_22), .down(vreg_20_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_21), .sw(sw));
	wire signed[17:0] vwire_20_22;
	reg signed[17:0] vreg_20_22;
	node n20_22(.left(vreg_19_22), .right(vreg_21_22), .up(vreg_20_23), .down(vreg_20_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_22), .sw(sw));
	wire signed[17:0] vwire_20_23;
	reg signed[17:0] vreg_20_23;
	node n20_23(.left(vreg_19_23), .right(vreg_21_23), .up(vreg_20_24), .down(vreg_20_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_23), .sw(sw));
	wire signed[17:0] vwire_20_24;
	reg signed[17:0] vreg_20_24;
	node n20_24(.left(vreg_19_24), .right(vreg_21_24), .up(vreg_20_25), .down(vreg_20_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_24), .sw(sw));
	wire signed[17:0] vwire_20_25;
	reg signed[17:0] vreg_20_25;
	node n20_25(.left(vreg_19_25), .right(vreg_21_25), .up(vreg_20_26), .down(vreg_20_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_25), .sw(sw));
	wire signed[17:0] vwire_20_26;
	reg signed[17:0] vreg_20_26;
	node n20_26(.left(vreg_19_26), .right(vreg_21_26), .up(vreg_20_27), .down(vreg_20_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_26), .sw(sw));
	wire signed[17:0] vwire_20_27;
	reg signed[17:0] vreg_20_27;
	node n20_27(.left(vreg_19_27), .right(vreg_21_27), .up(vreg_20_28), .down(vreg_20_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_27), .sw(sw));
	wire signed[17:0] vwire_20_28;
	reg signed[17:0] vreg_20_28;
	node n20_28(.left(vreg_19_28), .right(vreg_21_28), .up(vreg_20_29), .down(vreg_20_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_28), .sw(sw));
	wire signed[17:0] vwire_20_29;
	reg signed[17:0] vreg_20_29;
	node n20_29(.left(vreg_19_29), .right(vreg_21_29), .up(vreg_20_30), .down(vreg_20_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_29), .sw(sw));
	wire signed[17:0] vwire_20_30;
	reg signed[17:0] vreg_20_30;
	node n20_30(.left(vreg_19_30), .right(vreg_21_30), .up(vreg_20_31), .down(vreg_20_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_30), .sw(sw));
	wire signed[17:0] vwire_20_31;
	reg signed[17:0] vreg_20_31;
	node n20_31(.left(vreg_19_31), .right(vreg_21_31), .up(vreg_20_32), .down(vreg_20_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_31), .sw(sw));
	wire signed[17:0] vwire_20_32;
	reg signed[17:0] vreg_20_32;
	node n20_32(.left(vreg_19_32), .right(vreg_21_32), .up(vreg_20_33), .down(vreg_20_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_32), .sw(sw));
	wire signed[17:0] vwire_20_33;
	reg signed[17:0] vreg_20_33;
	node n20_33(.left(vreg_19_33), .right(vreg_21_33), .up(vreg_20_34), .down(vreg_20_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_33), .sw(sw));
	wire signed[17:0] vwire_20_34;
	reg signed[17:0] vreg_20_34;
	node n20_34(.left(vreg_19_34), .right(vreg_21_34), .up(vreg_20_35), .down(vreg_20_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_34), .sw(sw));
	wire signed[17:0] vwire_20_35;
	reg signed[17:0] vreg_20_35;
	node n20_35(.left(vreg_19_35), .right(vreg_21_35), .up(vreg_20_36), .down(vreg_20_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_35), .sw(sw));
	wire signed[17:0] vwire_20_36;
	reg signed[17:0] vreg_20_36;
	node n20_36(.left(vreg_19_36), .right(vreg_21_36), .up(vreg_20_37), .down(vreg_20_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_36), .sw(sw));
	wire signed[17:0] vwire_20_37;
	reg signed[17:0] vreg_20_37;
	node n20_37(.left(vreg_19_37), .right(vreg_21_37), .up(vreg_20_38), .down(vreg_20_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_37), .sw(sw));
	wire signed[17:0] vwire_20_38;
	reg signed[17:0] vreg_20_38;
	node n20_38(.left(vreg_19_38), .right(vreg_21_38), .up(vreg_20_39), .down(vreg_20_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_38), .sw(sw));
	wire signed[17:0] vwire_20_39;
	reg signed[17:0] vreg_20_39;
	node n20_39(.left(vreg_19_39), .right(vreg_21_39), .up(vreg_20_40), .down(vreg_20_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_39), .sw(sw));
	wire signed[17:0] vwire_20_40;
	reg signed[17:0] vreg_20_40;
	node n20_40(.left(vreg_19_40), .right(vreg_21_40), .up(vreg_20_41), .down(vreg_20_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_40), .sw(sw));
	wire signed[17:0] vwire_20_41;
	reg signed[17:0] vreg_20_41;
	node n20_41(.left(vreg_19_41), .right(vreg_21_41), .up(vreg_20_42), .down(vreg_20_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_41), .sw(sw));
	wire signed[17:0] vwire_20_42;
	reg signed[17:0] vreg_20_42;
	node n20_42(.left(vreg_19_42), .right(vreg_21_42), .up(vreg_20_43), .down(vreg_20_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_42), .sw(sw));
	wire signed[17:0] vwire_20_43;
	reg signed[17:0] vreg_20_43;
	node n20_43(.left(vreg_19_43), .right(vreg_21_43), .up(vreg_20_44), .down(vreg_20_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_43), .sw(sw));
	wire signed[17:0] vwire_20_44;
	reg signed[17:0] vreg_20_44;
	node n20_44(.left(vreg_19_44), .right(vreg_21_44), .up(vreg_20_45), .down(vreg_20_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_44), .sw(sw));
	wire signed[17:0] vwire_20_45;
	reg signed[17:0] vreg_20_45;
	node n20_45(.left(vreg_19_45), .right(vreg_21_45), .up(vreg_20_46), .down(vreg_20_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_45), .sw(sw));
	wire signed[17:0] vwire_20_46;
	reg signed[17:0] vreg_20_46;
	node n20_46(.left(vreg_19_46), .right(vreg_21_46), .up(vreg_20_47), .down(vreg_20_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_46), .sw(sw));
	wire signed[17:0] vwire_20_47;
	reg signed[17:0] vreg_20_47;
	node n20_47(.left(vreg_19_47), .right(vreg_21_47), .up(vreg_20_48), .down(vreg_20_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_47), .sw(sw));
	wire signed[17:0] vwire_20_48;
	reg signed[17:0] vreg_20_48;
	node n20_48(.left(vreg_19_48), .right(vreg_21_48), .up(vreg_20_49), .down(vreg_20_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_48), .sw(sw));
	wire signed[17:0] vwire_20_49;
	reg signed[17:0] vreg_20_49;
	node n20_49(.left(vreg_19_49), .right(vreg_21_49), .up(18'b0), .down(vreg_20_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_20_49), .sw(sw));
	wire signed[17:0] vwire_21_0;
	reg signed[17:0] vreg_21_0;
	node n21_0(.left(vreg_20_0), .right(vreg_22_0), .up(vreg_21_1), .down(vreg_21_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_0), .sw(sw));
	wire signed[17:0] vwire_21_1;
	reg signed[17:0] vreg_21_1;
	node n21_1(.left(vreg_20_1), .right(vreg_22_1), .up(vreg_21_2), .down(vreg_21_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_1), .sw(sw));
	wire signed[17:0] vwire_21_2;
	reg signed[17:0] vreg_21_2;
	node n21_2(.left(vreg_20_2), .right(vreg_22_2), .up(vreg_21_3), .down(vreg_21_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_2), .sw(sw));
	wire signed[17:0] vwire_21_3;
	reg signed[17:0] vreg_21_3;
	node n21_3(.left(vreg_20_3), .right(vreg_22_3), .up(vreg_21_4), .down(vreg_21_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_3), .sw(sw));
	wire signed[17:0] vwire_21_4;
	reg signed[17:0] vreg_21_4;
	node n21_4(.left(vreg_20_4), .right(vreg_22_4), .up(vreg_21_5), .down(vreg_21_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_4), .sw(sw));
	wire signed[17:0] vwire_21_5;
	reg signed[17:0] vreg_21_5;
	node n21_5(.left(vreg_20_5), .right(vreg_22_5), .up(vreg_21_6), .down(vreg_21_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_5), .sw(sw));
	wire signed[17:0] vwire_21_6;
	reg signed[17:0] vreg_21_6;
	node n21_6(.left(vreg_20_6), .right(vreg_22_6), .up(vreg_21_7), .down(vreg_21_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_6), .sw(sw));
	wire signed[17:0] vwire_21_7;
	reg signed[17:0] vreg_21_7;
	node n21_7(.left(vreg_20_7), .right(vreg_22_7), .up(vreg_21_8), .down(vreg_21_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_7), .sw(sw));
	wire signed[17:0] vwire_21_8;
	reg signed[17:0] vreg_21_8;
	node n21_8(.left(vreg_20_8), .right(vreg_22_8), .up(vreg_21_9), .down(vreg_21_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_8), .sw(sw));
	wire signed[17:0] vwire_21_9;
	reg signed[17:0] vreg_21_9;
	node n21_9(.left(vreg_20_9), .right(vreg_22_9), .up(vreg_21_10), .down(vreg_21_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_9), .sw(sw));
	wire signed[17:0] vwire_21_10;
	reg signed[17:0] vreg_21_10;
	node n21_10(.left(vreg_20_10), .right(vreg_22_10), .up(vreg_21_11), .down(vreg_21_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_10), .sw(sw));
	wire signed[17:0] vwire_21_11;
	reg signed[17:0] vreg_21_11;
	node n21_11(.left(vreg_20_11), .right(vreg_22_11), .up(vreg_21_12), .down(vreg_21_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_11), .sw(sw));
	wire signed[17:0] vwire_21_12;
	reg signed[17:0] vreg_21_12;
	node n21_12(.left(vreg_20_12), .right(vreg_22_12), .up(vreg_21_13), .down(vreg_21_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_12), .sw(sw));
	wire signed[17:0] vwire_21_13;
	reg signed[17:0] vreg_21_13;
	node n21_13(.left(vreg_20_13), .right(vreg_22_13), .up(vreg_21_14), .down(vreg_21_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_13), .sw(sw));
	wire signed[17:0] vwire_21_14;
	reg signed[17:0] vreg_21_14;
	node n21_14(.left(vreg_20_14), .right(vreg_22_14), .up(vreg_21_15), .down(vreg_21_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_14), .sw(sw));
	wire signed[17:0] vwire_21_15;
	reg signed[17:0] vreg_21_15;
	node n21_15(.left(vreg_20_15), .right(vreg_22_15), .up(vreg_21_16), .down(vreg_21_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_15), .sw(sw));
	wire signed[17:0] vwire_21_16;
	reg signed[17:0] vreg_21_16;
	node n21_16(.left(vreg_20_16), .right(vreg_22_16), .up(vreg_21_17), .down(vreg_21_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_16), .sw(sw));
	wire signed[17:0] vwire_21_17;
	reg signed[17:0] vreg_21_17;
	node n21_17(.left(vreg_20_17), .right(vreg_22_17), .up(vreg_21_18), .down(vreg_21_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_17), .sw(sw));
	wire signed[17:0] vwire_21_18;
	reg signed[17:0] vreg_21_18;
	node n21_18(.left(vreg_20_18), .right(vreg_22_18), .up(vreg_21_19), .down(vreg_21_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_18), .sw(sw));
	wire signed[17:0] vwire_21_19;
	reg signed[17:0] vreg_21_19;
	node n21_19(.left(vreg_20_19), .right(vreg_22_19), .up(vreg_21_20), .down(vreg_21_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_19), .sw(sw));
	wire signed[17:0] vwire_21_20;
	reg signed[17:0] vreg_21_20;
	node n21_20(.left(vreg_20_20), .right(vreg_22_20), .up(vreg_21_21), .down(vreg_21_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_20), .sw(sw));
	wire signed[17:0] vwire_21_21;
	reg signed[17:0] vreg_21_21;
	node n21_21(.left(vreg_20_21), .right(vreg_22_21), .up(vreg_21_22), .down(vreg_21_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_21), .sw(sw));
	wire signed[17:0] vwire_21_22;
	reg signed[17:0] vreg_21_22;
	node n21_22(.left(vreg_20_22), .right(vreg_22_22), .up(vreg_21_23), .down(vreg_21_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_22), .sw(sw));
	wire signed[17:0] vwire_21_23;
	reg signed[17:0] vreg_21_23;
	node n21_23(.left(vreg_20_23), .right(vreg_22_23), .up(vreg_21_24), .down(vreg_21_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_23), .sw(sw));
	wire signed[17:0] vwire_21_24;
	reg signed[17:0] vreg_21_24;
	node n21_24(.left(vreg_20_24), .right(vreg_22_24), .up(vreg_21_25), .down(vreg_21_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_24), .sw(sw));
	wire signed[17:0] vwire_21_25;
	reg signed[17:0] vreg_21_25;
	node n21_25(.left(vreg_20_25), .right(vreg_22_25), .up(vreg_21_26), .down(vreg_21_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_25), .sw(sw));
	wire signed[17:0] vwire_21_26;
	reg signed[17:0] vreg_21_26;
	node n21_26(.left(vreg_20_26), .right(vreg_22_26), .up(vreg_21_27), .down(vreg_21_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_26), .sw(sw));
	wire signed[17:0] vwire_21_27;
	reg signed[17:0] vreg_21_27;
	node n21_27(.left(vreg_20_27), .right(vreg_22_27), .up(vreg_21_28), .down(vreg_21_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_27), .sw(sw));
	wire signed[17:0] vwire_21_28;
	reg signed[17:0] vreg_21_28;
	node n21_28(.left(vreg_20_28), .right(vreg_22_28), .up(vreg_21_29), .down(vreg_21_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_28), .sw(sw));
	wire signed[17:0] vwire_21_29;
	reg signed[17:0] vreg_21_29;
	node n21_29(.left(vreg_20_29), .right(vreg_22_29), .up(vreg_21_30), .down(vreg_21_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_29), .sw(sw));
	wire signed[17:0] vwire_21_30;
	reg signed[17:0] vreg_21_30;
	node n21_30(.left(vreg_20_30), .right(vreg_22_30), .up(vreg_21_31), .down(vreg_21_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_30), .sw(sw));
	wire signed[17:0] vwire_21_31;
	reg signed[17:0] vreg_21_31;
	node n21_31(.left(vreg_20_31), .right(vreg_22_31), .up(vreg_21_32), .down(vreg_21_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_31), .sw(sw));
	wire signed[17:0] vwire_21_32;
	reg signed[17:0] vreg_21_32;
	node n21_32(.left(vreg_20_32), .right(vreg_22_32), .up(vreg_21_33), .down(vreg_21_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_32), .sw(sw));
	wire signed[17:0] vwire_21_33;
	reg signed[17:0] vreg_21_33;
	node n21_33(.left(vreg_20_33), .right(vreg_22_33), .up(vreg_21_34), .down(vreg_21_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_33), .sw(sw));
	wire signed[17:0] vwire_21_34;
	reg signed[17:0] vreg_21_34;
	node n21_34(.left(vreg_20_34), .right(vreg_22_34), .up(vreg_21_35), .down(vreg_21_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_34), .sw(sw));
	wire signed[17:0] vwire_21_35;
	reg signed[17:0] vreg_21_35;
	node n21_35(.left(vreg_20_35), .right(vreg_22_35), .up(vreg_21_36), .down(vreg_21_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_35), .sw(sw));
	wire signed[17:0] vwire_21_36;
	reg signed[17:0] vreg_21_36;
	node n21_36(.left(vreg_20_36), .right(vreg_22_36), .up(vreg_21_37), .down(vreg_21_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_36), .sw(sw));
	wire signed[17:0] vwire_21_37;
	reg signed[17:0] vreg_21_37;
	node n21_37(.left(vreg_20_37), .right(vreg_22_37), .up(vreg_21_38), .down(vreg_21_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_37), .sw(sw));
	wire signed[17:0] vwire_21_38;
	reg signed[17:0] vreg_21_38;
	node n21_38(.left(vreg_20_38), .right(vreg_22_38), .up(vreg_21_39), .down(vreg_21_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_38), .sw(sw));
	wire signed[17:0] vwire_21_39;
	reg signed[17:0] vreg_21_39;
	node n21_39(.left(vreg_20_39), .right(vreg_22_39), .up(vreg_21_40), .down(vreg_21_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_39), .sw(sw));
	wire signed[17:0] vwire_21_40;
	reg signed[17:0] vreg_21_40;
	node n21_40(.left(vreg_20_40), .right(vreg_22_40), .up(vreg_21_41), .down(vreg_21_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_40), .sw(sw));
	wire signed[17:0] vwire_21_41;
	reg signed[17:0] vreg_21_41;
	node n21_41(.left(vreg_20_41), .right(vreg_22_41), .up(vreg_21_42), .down(vreg_21_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_41), .sw(sw));
	wire signed[17:0] vwire_21_42;
	reg signed[17:0] vreg_21_42;
	node n21_42(.left(vreg_20_42), .right(vreg_22_42), .up(vreg_21_43), .down(vreg_21_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_42), .sw(sw));
	wire signed[17:0] vwire_21_43;
	reg signed[17:0] vreg_21_43;
	node n21_43(.left(vreg_20_43), .right(vreg_22_43), .up(vreg_21_44), .down(vreg_21_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_43), .sw(sw));
	wire signed[17:0] vwire_21_44;
	reg signed[17:0] vreg_21_44;
	node n21_44(.left(vreg_20_44), .right(vreg_22_44), .up(vreg_21_45), .down(vreg_21_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_44), .sw(sw));
	wire signed[17:0] vwire_21_45;
	reg signed[17:0] vreg_21_45;
	node n21_45(.left(vreg_20_45), .right(vreg_22_45), .up(vreg_21_46), .down(vreg_21_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_45), .sw(sw));
	wire signed[17:0] vwire_21_46;
	reg signed[17:0] vreg_21_46;
	node n21_46(.left(vreg_20_46), .right(vreg_22_46), .up(vreg_21_47), .down(vreg_21_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_46), .sw(sw));
	wire signed[17:0] vwire_21_47;
	reg signed[17:0] vreg_21_47;
	node n21_47(.left(vreg_20_47), .right(vreg_22_47), .up(vreg_21_48), .down(vreg_21_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_47), .sw(sw));
	wire signed[17:0] vwire_21_48;
	reg signed[17:0] vreg_21_48;
	node n21_48(.left(vreg_20_48), .right(vreg_22_48), .up(vreg_21_49), .down(vreg_21_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_48), .sw(sw));
	wire signed[17:0] vwire_21_49;
	reg signed[17:0] vreg_21_49;
	node n21_49(.left(vreg_20_49), .right(vreg_22_49), .up(18'b0), .down(vreg_21_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_21_49), .sw(sw));
	wire signed[17:0] vwire_22_0;
	reg signed[17:0] vreg_22_0;
	node n22_0(.left(vreg_21_0), .right(vreg_23_0), .up(vreg_22_1), .down(vreg_22_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_0), .sw(sw));
	wire signed[17:0] vwire_22_1;
	reg signed[17:0] vreg_22_1;
	node n22_1(.left(vreg_21_1), .right(vreg_23_1), .up(vreg_22_2), .down(vreg_22_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_1), .sw(sw));
	wire signed[17:0] vwire_22_2;
	reg signed[17:0] vreg_22_2;
	node n22_2(.left(vreg_21_2), .right(vreg_23_2), .up(vreg_22_3), .down(vreg_22_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_2), .sw(sw));
	wire signed[17:0] vwire_22_3;
	reg signed[17:0] vreg_22_3;
	node n22_3(.left(vreg_21_3), .right(vreg_23_3), .up(vreg_22_4), .down(vreg_22_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_3), .sw(sw));
	wire signed[17:0] vwire_22_4;
	reg signed[17:0] vreg_22_4;
	node n22_4(.left(vreg_21_4), .right(vreg_23_4), .up(vreg_22_5), .down(vreg_22_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_4), .sw(sw));
	wire signed[17:0] vwire_22_5;
	reg signed[17:0] vreg_22_5;
	node n22_5(.left(vreg_21_5), .right(vreg_23_5), .up(vreg_22_6), .down(vreg_22_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_5), .sw(sw));
	wire signed[17:0] vwire_22_6;
	reg signed[17:0] vreg_22_6;
	node n22_6(.left(vreg_21_6), .right(vreg_23_6), .up(vreg_22_7), .down(vreg_22_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_6), .sw(sw));
	wire signed[17:0] vwire_22_7;
	reg signed[17:0] vreg_22_7;
	node n22_7(.left(vreg_21_7), .right(vreg_23_7), .up(vreg_22_8), .down(vreg_22_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_7), .sw(sw));
	wire signed[17:0] vwire_22_8;
	reg signed[17:0] vreg_22_8;
	node n22_8(.left(vreg_21_8), .right(vreg_23_8), .up(vreg_22_9), .down(vreg_22_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_8), .sw(sw));
	wire signed[17:0] vwire_22_9;
	reg signed[17:0] vreg_22_9;
	node n22_9(.left(vreg_21_9), .right(vreg_23_9), .up(vreg_22_10), .down(vreg_22_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_9), .sw(sw));
	wire signed[17:0] vwire_22_10;
	reg signed[17:0] vreg_22_10;
	node n22_10(.left(vreg_21_10), .right(vreg_23_10), .up(vreg_22_11), .down(vreg_22_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_10), .sw(sw));
	wire signed[17:0] vwire_22_11;
	reg signed[17:0] vreg_22_11;
	node n22_11(.left(vreg_21_11), .right(vreg_23_11), .up(vreg_22_12), .down(vreg_22_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_11), .sw(sw));
	wire signed[17:0] vwire_22_12;
	reg signed[17:0] vreg_22_12;
	node n22_12(.left(vreg_21_12), .right(vreg_23_12), .up(vreg_22_13), .down(vreg_22_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_12), .sw(sw));
	wire signed[17:0] vwire_22_13;
	reg signed[17:0] vreg_22_13;
	node n22_13(.left(vreg_21_13), .right(vreg_23_13), .up(vreg_22_14), .down(vreg_22_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_13), .sw(sw));
	wire signed[17:0] vwire_22_14;
	reg signed[17:0] vreg_22_14;
	node n22_14(.left(vreg_21_14), .right(vreg_23_14), .up(vreg_22_15), .down(vreg_22_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_14), .sw(sw));
	wire signed[17:0] vwire_22_15;
	reg signed[17:0] vreg_22_15;
	node n22_15(.left(vreg_21_15), .right(vreg_23_15), .up(vreg_22_16), .down(vreg_22_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_15), .sw(sw));
	wire signed[17:0] vwire_22_16;
	reg signed[17:0] vreg_22_16;
	node n22_16(.left(vreg_21_16), .right(vreg_23_16), .up(vreg_22_17), .down(vreg_22_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_16), .sw(sw));
	wire signed[17:0] vwire_22_17;
	reg signed[17:0] vreg_22_17;
	node n22_17(.left(vreg_21_17), .right(vreg_23_17), .up(vreg_22_18), .down(vreg_22_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_17), .sw(sw));
	wire signed[17:0] vwire_22_18;
	reg signed[17:0] vreg_22_18;
	node n22_18(.left(vreg_21_18), .right(vreg_23_18), .up(vreg_22_19), .down(vreg_22_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_18), .sw(sw));
	wire signed[17:0] vwire_22_19;
	reg signed[17:0] vreg_22_19;
	node n22_19(.left(vreg_21_19), .right(vreg_23_19), .up(vreg_22_20), .down(vreg_22_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_19), .sw(sw));
	wire signed[17:0] vwire_22_20;
	reg signed[17:0] vreg_22_20;
	node n22_20(.left(vreg_21_20), .right(vreg_23_20), .up(vreg_22_21), .down(vreg_22_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_20), .sw(sw));
	wire signed[17:0] vwire_22_21;
	reg signed[17:0] vreg_22_21;
	node n22_21(.left(vreg_21_21), .right(vreg_23_21), .up(vreg_22_22), .down(vreg_22_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_21), .sw(sw));
	wire signed[17:0] vwire_22_22;
	reg signed[17:0] vreg_22_22;
	node n22_22(.left(vreg_21_22), .right(vreg_23_22), .up(vreg_22_23), .down(vreg_22_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_22), .sw(sw));
	wire signed[17:0] vwire_22_23;
	reg signed[17:0] vreg_22_23;
	node n22_23(.left(vreg_21_23), .right(vreg_23_23), .up(vreg_22_24), .down(vreg_22_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_23), .sw(sw));
	wire signed[17:0] vwire_22_24;
	reg signed[17:0] vreg_22_24;
	node n22_24(.left(vreg_21_24), .right(vreg_23_24), .up(vreg_22_25), .down(vreg_22_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_24), .sw(sw));
	wire signed[17:0] vwire_22_25;
	reg signed[17:0] vreg_22_25;
	node n22_25(.left(vreg_21_25), .right(vreg_23_25), .up(vreg_22_26), .down(vreg_22_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_25), .sw(sw));
	wire signed[17:0] vwire_22_26;
	reg signed[17:0] vreg_22_26;
	node n22_26(.left(vreg_21_26), .right(vreg_23_26), .up(vreg_22_27), .down(vreg_22_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_26), .sw(sw));
	wire signed[17:0] vwire_22_27;
	reg signed[17:0] vreg_22_27;
	node n22_27(.left(vreg_21_27), .right(vreg_23_27), .up(vreg_22_28), .down(vreg_22_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_27), .sw(sw));
	wire signed[17:0] vwire_22_28;
	reg signed[17:0] vreg_22_28;
	node n22_28(.left(vreg_21_28), .right(vreg_23_28), .up(vreg_22_29), .down(vreg_22_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_28), .sw(sw));
	wire signed[17:0] vwire_22_29;
	reg signed[17:0] vreg_22_29;
	node n22_29(.left(vreg_21_29), .right(vreg_23_29), .up(vreg_22_30), .down(vreg_22_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_29), .sw(sw));
	wire signed[17:0] vwire_22_30;
	reg signed[17:0] vreg_22_30;
	node n22_30(.left(vreg_21_30), .right(vreg_23_30), .up(vreg_22_31), .down(vreg_22_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_30), .sw(sw));
	wire signed[17:0] vwire_22_31;
	reg signed[17:0] vreg_22_31;
	node n22_31(.left(vreg_21_31), .right(vreg_23_31), .up(vreg_22_32), .down(vreg_22_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_31), .sw(sw));
	wire signed[17:0] vwire_22_32;
	reg signed[17:0] vreg_22_32;
	node n22_32(.left(vreg_21_32), .right(vreg_23_32), .up(vreg_22_33), .down(vreg_22_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_32), .sw(sw));
	wire signed[17:0] vwire_22_33;
	reg signed[17:0] vreg_22_33;
	node n22_33(.left(vreg_21_33), .right(vreg_23_33), .up(vreg_22_34), .down(vreg_22_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_33), .sw(sw));
	wire signed[17:0] vwire_22_34;
	reg signed[17:0] vreg_22_34;
	node n22_34(.left(vreg_21_34), .right(vreg_23_34), .up(vreg_22_35), .down(vreg_22_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_34), .sw(sw));
	wire signed[17:0] vwire_22_35;
	reg signed[17:0] vreg_22_35;
	node n22_35(.left(vreg_21_35), .right(vreg_23_35), .up(vreg_22_36), .down(vreg_22_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_35), .sw(sw));
	wire signed[17:0] vwire_22_36;
	reg signed[17:0] vreg_22_36;
	node n22_36(.left(vreg_21_36), .right(vreg_23_36), .up(vreg_22_37), .down(vreg_22_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_36), .sw(sw));
	wire signed[17:0] vwire_22_37;
	reg signed[17:0] vreg_22_37;
	node n22_37(.left(vreg_21_37), .right(vreg_23_37), .up(vreg_22_38), .down(vreg_22_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_37), .sw(sw));
	wire signed[17:0] vwire_22_38;
	reg signed[17:0] vreg_22_38;
	node n22_38(.left(vreg_21_38), .right(vreg_23_38), .up(vreg_22_39), .down(vreg_22_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_38), .sw(sw));
	wire signed[17:0] vwire_22_39;
	reg signed[17:0] vreg_22_39;
	node n22_39(.left(vreg_21_39), .right(vreg_23_39), .up(vreg_22_40), .down(vreg_22_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_39), .sw(sw));
	wire signed[17:0] vwire_22_40;
	reg signed[17:0] vreg_22_40;
	node n22_40(.left(vreg_21_40), .right(vreg_23_40), .up(vreg_22_41), .down(vreg_22_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_40), .sw(sw));
	wire signed[17:0] vwire_22_41;
	reg signed[17:0] vreg_22_41;
	node n22_41(.left(vreg_21_41), .right(vreg_23_41), .up(vreg_22_42), .down(vreg_22_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_41), .sw(sw));
	wire signed[17:0] vwire_22_42;
	reg signed[17:0] vreg_22_42;
	node n22_42(.left(vreg_21_42), .right(vreg_23_42), .up(vreg_22_43), .down(vreg_22_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_42), .sw(sw));
	wire signed[17:0] vwire_22_43;
	reg signed[17:0] vreg_22_43;
	node n22_43(.left(vreg_21_43), .right(vreg_23_43), .up(vreg_22_44), .down(vreg_22_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_43), .sw(sw));
	wire signed[17:0] vwire_22_44;
	reg signed[17:0] vreg_22_44;
	node n22_44(.left(vreg_21_44), .right(vreg_23_44), .up(vreg_22_45), .down(vreg_22_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_44), .sw(sw));
	wire signed[17:0] vwire_22_45;
	reg signed[17:0] vreg_22_45;
	node n22_45(.left(vreg_21_45), .right(vreg_23_45), .up(vreg_22_46), .down(vreg_22_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_45), .sw(sw));
	wire signed[17:0] vwire_22_46;
	reg signed[17:0] vreg_22_46;
	node n22_46(.left(vreg_21_46), .right(vreg_23_46), .up(vreg_22_47), .down(vreg_22_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_46), .sw(sw));
	wire signed[17:0] vwire_22_47;
	reg signed[17:0] vreg_22_47;
	node n22_47(.left(vreg_21_47), .right(vreg_23_47), .up(vreg_22_48), .down(vreg_22_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_47), .sw(sw));
	wire signed[17:0] vwire_22_48;
	reg signed[17:0] vreg_22_48;
	node n22_48(.left(vreg_21_48), .right(vreg_23_48), .up(vreg_22_49), .down(vreg_22_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_48), .sw(sw));
	wire signed[17:0] vwire_22_49;
	reg signed[17:0] vreg_22_49;
	node n22_49(.left(vreg_21_49), .right(vreg_23_49), .up(18'b0), .down(vreg_22_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_22_49), .sw(sw));
	wire signed[17:0] vwire_23_0;
	reg signed[17:0] vreg_23_0;
	node n23_0(.left(vreg_22_0), .right(vreg_24_0), .up(vreg_23_1), .down(vreg_23_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_0), .sw(sw));
	wire signed[17:0] vwire_23_1;
	reg signed[17:0] vreg_23_1;
	node n23_1(.left(vreg_22_1), .right(vreg_24_1), .up(vreg_23_2), .down(vreg_23_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_1), .sw(sw));
	wire signed[17:0] vwire_23_2;
	reg signed[17:0] vreg_23_2;
	node n23_2(.left(vreg_22_2), .right(vreg_24_2), .up(vreg_23_3), .down(vreg_23_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_2), .sw(sw));
	wire signed[17:0] vwire_23_3;
	reg signed[17:0] vreg_23_3;
	node n23_3(.left(vreg_22_3), .right(vreg_24_3), .up(vreg_23_4), .down(vreg_23_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_3), .sw(sw));
	wire signed[17:0] vwire_23_4;
	reg signed[17:0] vreg_23_4;
	node n23_4(.left(vreg_22_4), .right(vreg_24_4), .up(vreg_23_5), .down(vreg_23_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_4), .sw(sw));
	wire signed[17:0] vwire_23_5;
	reg signed[17:0] vreg_23_5;
	node n23_5(.left(vreg_22_5), .right(vreg_24_5), .up(vreg_23_6), .down(vreg_23_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_5), .sw(sw));
	wire signed[17:0] vwire_23_6;
	reg signed[17:0] vreg_23_6;
	node n23_6(.left(vreg_22_6), .right(vreg_24_6), .up(vreg_23_7), .down(vreg_23_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_6), .sw(sw));
	wire signed[17:0] vwire_23_7;
	reg signed[17:0] vreg_23_7;
	node n23_7(.left(vreg_22_7), .right(vreg_24_7), .up(vreg_23_8), .down(vreg_23_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_7), .sw(sw));
	wire signed[17:0] vwire_23_8;
	reg signed[17:0] vreg_23_8;
	node n23_8(.left(vreg_22_8), .right(vreg_24_8), .up(vreg_23_9), .down(vreg_23_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_8), .sw(sw));
	wire signed[17:0] vwire_23_9;
	reg signed[17:0] vreg_23_9;
	node n23_9(.left(vreg_22_9), .right(vreg_24_9), .up(vreg_23_10), .down(vreg_23_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_9), .sw(sw));
	wire signed[17:0] vwire_23_10;
	reg signed[17:0] vreg_23_10;
	node n23_10(.left(vreg_22_10), .right(vreg_24_10), .up(vreg_23_11), .down(vreg_23_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_10), .sw(sw));
	wire signed[17:0] vwire_23_11;
	reg signed[17:0] vreg_23_11;
	node n23_11(.left(vreg_22_11), .right(vreg_24_11), .up(vreg_23_12), .down(vreg_23_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_11), .sw(sw));
	wire signed[17:0] vwire_23_12;
	reg signed[17:0] vreg_23_12;
	node n23_12(.left(vreg_22_12), .right(vreg_24_12), .up(vreg_23_13), .down(vreg_23_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_12), .sw(sw));
	wire signed[17:0] vwire_23_13;
	reg signed[17:0] vreg_23_13;
	node n23_13(.left(vreg_22_13), .right(vreg_24_13), .up(vreg_23_14), .down(vreg_23_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_13), .sw(sw));
	wire signed[17:0] vwire_23_14;
	reg signed[17:0] vreg_23_14;
	node n23_14(.left(vreg_22_14), .right(vreg_24_14), .up(vreg_23_15), .down(vreg_23_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_14), .sw(sw));
	wire signed[17:0] vwire_23_15;
	reg signed[17:0] vreg_23_15;
	node n23_15(.left(vreg_22_15), .right(vreg_24_15), .up(vreg_23_16), .down(vreg_23_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_15), .sw(sw));
	wire signed[17:0] vwire_23_16;
	reg signed[17:0] vreg_23_16;
	node n23_16(.left(vreg_22_16), .right(vreg_24_16), .up(vreg_23_17), .down(vreg_23_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_16), .sw(sw));
	wire signed[17:0] vwire_23_17;
	reg signed[17:0] vreg_23_17;
	node n23_17(.left(vreg_22_17), .right(vreg_24_17), .up(vreg_23_18), .down(vreg_23_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_17), .sw(sw));
	wire signed[17:0] vwire_23_18;
	reg signed[17:0] vreg_23_18;
	node n23_18(.left(vreg_22_18), .right(vreg_24_18), .up(vreg_23_19), .down(vreg_23_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_18), .sw(sw));
	wire signed[17:0] vwire_23_19;
	reg signed[17:0] vreg_23_19;
	node n23_19(.left(vreg_22_19), .right(vreg_24_19), .up(vreg_23_20), .down(vreg_23_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_19), .sw(sw));
	wire signed[17:0] vwire_23_20;
	reg signed[17:0] vreg_23_20;
	node n23_20(.left(vreg_22_20), .right(vreg_24_20), .up(vreg_23_21), .down(vreg_23_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_20), .sw(sw));
	wire signed[17:0] vwire_23_21;
	reg signed[17:0] vreg_23_21;
	node n23_21(.left(vreg_22_21), .right(vreg_24_21), .up(vreg_23_22), .down(vreg_23_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_21), .sw(sw));
	wire signed[17:0] vwire_23_22;
	reg signed[17:0] vreg_23_22;
	node n23_22(.left(vreg_22_22), .right(vreg_24_22), .up(vreg_23_23), .down(vreg_23_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_22), .sw(sw));
	wire signed[17:0] vwire_23_23;
	reg signed[17:0] vreg_23_23;
	node n23_23(.left(vreg_22_23), .right(vreg_24_23), .up(vreg_23_24), .down(vreg_23_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_23), .sw(sw));
	wire signed[17:0] vwire_23_24;
	reg signed[17:0] vreg_23_24;
	node n23_24(.left(vreg_22_24), .right(vreg_24_24), .up(vreg_23_25), .down(vreg_23_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_24), .sw(sw));
	wire signed[17:0] vwire_23_25;
	reg signed[17:0] vreg_23_25;
	node n23_25(.left(vreg_22_25), .right(vreg_24_25), .up(vreg_23_26), .down(vreg_23_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_25), .sw(sw));
	wire signed[17:0] vwire_23_26;
	reg signed[17:0] vreg_23_26;
	node n23_26(.left(vreg_22_26), .right(vreg_24_26), .up(vreg_23_27), .down(vreg_23_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_26), .sw(sw));
	wire signed[17:0] vwire_23_27;
	reg signed[17:0] vreg_23_27;
	node n23_27(.left(vreg_22_27), .right(vreg_24_27), .up(vreg_23_28), .down(vreg_23_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_27), .sw(sw));
	wire signed[17:0] vwire_23_28;
	reg signed[17:0] vreg_23_28;
	node n23_28(.left(vreg_22_28), .right(vreg_24_28), .up(vreg_23_29), .down(vreg_23_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_28), .sw(sw));
	wire signed[17:0] vwire_23_29;
	reg signed[17:0] vreg_23_29;
	node n23_29(.left(vreg_22_29), .right(vreg_24_29), .up(vreg_23_30), .down(vreg_23_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_29), .sw(sw));
	wire signed[17:0] vwire_23_30;
	reg signed[17:0] vreg_23_30;
	node n23_30(.left(vreg_22_30), .right(vreg_24_30), .up(vreg_23_31), .down(vreg_23_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_30), .sw(sw));
	wire signed[17:0] vwire_23_31;
	reg signed[17:0] vreg_23_31;
	node n23_31(.left(vreg_22_31), .right(vreg_24_31), .up(vreg_23_32), .down(vreg_23_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_31), .sw(sw));
	wire signed[17:0] vwire_23_32;
	reg signed[17:0] vreg_23_32;
	node n23_32(.left(vreg_22_32), .right(vreg_24_32), .up(vreg_23_33), .down(vreg_23_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_32), .sw(sw));
	wire signed[17:0] vwire_23_33;
	reg signed[17:0] vreg_23_33;
	node n23_33(.left(vreg_22_33), .right(vreg_24_33), .up(vreg_23_34), .down(vreg_23_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_33), .sw(sw));
	wire signed[17:0] vwire_23_34;
	reg signed[17:0] vreg_23_34;
	node n23_34(.left(vreg_22_34), .right(vreg_24_34), .up(vreg_23_35), .down(vreg_23_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_34), .sw(sw));
	wire signed[17:0] vwire_23_35;
	reg signed[17:0] vreg_23_35;
	node n23_35(.left(vreg_22_35), .right(vreg_24_35), .up(vreg_23_36), .down(vreg_23_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_35), .sw(sw));
	wire signed[17:0] vwire_23_36;
	reg signed[17:0] vreg_23_36;
	node n23_36(.left(vreg_22_36), .right(vreg_24_36), .up(vreg_23_37), .down(vreg_23_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_36), .sw(sw));
	wire signed[17:0] vwire_23_37;
	reg signed[17:0] vreg_23_37;
	node n23_37(.left(vreg_22_37), .right(vreg_24_37), .up(vreg_23_38), .down(vreg_23_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_37), .sw(sw));
	wire signed[17:0] vwire_23_38;
	reg signed[17:0] vreg_23_38;
	node n23_38(.left(vreg_22_38), .right(vreg_24_38), .up(vreg_23_39), .down(vreg_23_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_38), .sw(sw));
	wire signed[17:0] vwire_23_39;
	reg signed[17:0] vreg_23_39;
	node n23_39(.left(vreg_22_39), .right(vreg_24_39), .up(vreg_23_40), .down(vreg_23_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_39), .sw(sw));
	wire signed[17:0] vwire_23_40;
	reg signed[17:0] vreg_23_40;
	node n23_40(.left(vreg_22_40), .right(vreg_24_40), .up(vreg_23_41), .down(vreg_23_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_40), .sw(sw));
	wire signed[17:0] vwire_23_41;
	reg signed[17:0] vreg_23_41;
	node n23_41(.left(vreg_22_41), .right(vreg_24_41), .up(vreg_23_42), .down(vreg_23_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_41), .sw(sw));
	wire signed[17:0] vwire_23_42;
	reg signed[17:0] vreg_23_42;
	node n23_42(.left(vreg_22_42), .right(vreg_24_42), .up(vreg_23_43), .down(vreg_23_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_42), .sw(sw));
	wire signed[17:0] vwire_23_43;
	reg signed[17:0] vreg_23_43;
	node n23_43(.left(vreg_22_43), .right(vreg_24_43), .up(vreg_23_44), .down(vreg_23_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_43), .sw(sw));
	wire signed[17:0] vwire_23_44;
	reg signed[17:0] vreg_23_44;
	node n23_44(.left(vreg_22_44), .right(vreg_24_44), .up(vreg_23_45), .down(vreg_23_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_44), .sw(sw));
	wire signed[17:0] vwire_23_45;
	reg signed[17:0] vreg_23_45;
	node n23_45(.left(vreg_22_45), .right(vreg_24_45), .up(vreg_23_46), .down(vreg_23_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_45), .sw(sw));
	wire signed[17:0] vwire_23_46;
	reg signed[17:0] vreg_23_46;
	node n23_46(.left(vreg_22_46), .right(vreg_24_46), .up(vreg_23_47), .down(vreg_23_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_46), .sw(sw));
	wire signed[17:0] vwire_23_47;
	reg signed[17:0] vreg_23_47;
	node n23_47(.left(vreg_22_47), .right(vreg_24_47), .up(vreg_23_48), .down(vreg_23_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_47), .sw(sw));
	wire signed[17:0] vwire_23_48;
	reg signed[17:0] vreg_23_48;
	node n23_48(.left(vreg_22_48), .right(vreg_24_48), .up(vreg_23_49), .down(vreg_23_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_48), .sw(sw));
	wire signed[17:0] vwire_23_49;
	reg signed[17:0] vreg_23_49;
	node n23_49(.left(vreg_22_49), .right(vreg_24_49), .up(18'b0), .down(vreg_23_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_23_49), .sw(sw));
	wire signed[17:0] vwire_24_0;
	reg signed[17:0] vreg_24_0;
	node n24_0(.left(vreg_23_0), .right(vreg_25_0), .up(vreg_24_1), .down(vreg_24_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_0), .sw(sw));
	wire signed[17:0] vwire_24_1;
	reg signed[17:0] vreg_24_1;
	node n24_1(.left(vreg_23_1), .right(vreg_25_1), .up(vreg_24_2), .down(vreg_24_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_1), .sw(sw));
	wire signed[17:0] vwire_24_2;
	reg signed[17:0] vreg_24_2;
	node n24_2(.left(vreg_23_2), .right(vreg_25_2), .up(vreg_24_3), .down(vreg_24_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_2), .sw(sw));
	wire signed[17:0] vwire_24_3;
	reg signed[17:0] vreg_24_3;
	node n24_3(.left(vreg_23_3), .right(vreg_25_3), .up(vreg_24_4), .down(vreg_24_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_3), .sw(sw));
	wire signed[17:0] vwire_24_4;
	reg signed[17:0] vreg_24_4;
	node n24_4(.left(vreg_23_4), .right(vreg_25_4), .up(vreg_24_5), .down(vreg_24_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_4), .sw(sw));
	wire signed[17:0] vwire_24_5;
	reg signed[17:0] vreg_24_5;
	node n24_5(.left(vreg_23_5), .right(vreg_25_5), .up(vreg_24_6), .down(vreg_24_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_5), .sw(sw));
	wire signed[17:0] vwire_24_6;
	reg signed[17:0] vreg_24_6;
	node n24_6(.left(vreg_23_6), .right(vreg_25_6), .up(vreg_24_7), .down(vreg_24_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_6), .sw(sw));
	wire signed[17:0] vwire_24_7;
	reg signed[17:0] vreg_24_7;
	node n24_7(.left(vreg_23_7), .right(vreg_25_7), .up(vreg_24_8), .down(vreg_24_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_7), .sw(sw));
	wire signed[17:0] vwire_24_8;
	reg signed[17:0] vreg_24_8;
	node n24_8(.left(vreg_23_8), .right(vreg_25_8), .up(vreg_24_9), .down(vreg_24_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_8), .sw(sw));
	wire signed[17:0] vwire_24_9;
	reg signed[17:0] vreg_24_9;
	node n24_9(.left(vreg_23_9), .right(vreg_25_9), .up(vreg_24_10), .down(vreg_24_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_9), .sw(sw));
	wire signed[17:0] vwire_24_10;
	reg signed[17:0] vreg_24_10;
	node n24_10(.left(vreg_23_10), .right(vreg_25_10), .up(vreg_24_11), .down(vreg_24_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_10), .sw(sw));
	wire signed[17:0] vwire_24_11;
	reg signed[17:0] vreg_24_11;
	node n24_11(.left(vreg_23_11), .right(vreg_25_11), .up(vreg_24_12), .down(vreg_24_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_11), .sw(sw));
	wire signed[17:0] vwire_24_12;
	reg signed[17:0] vreg_24_12;
	node n24_12(.left(vreg_23_12), .right(vreg_25_12), .up(vreg_24_13), .down(vreg_24_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_12), .sw(sw));
	wire signed[17:0] vwire_24_13;
	reg signed[17:0] vreg_24_13;
	node n24_13(.left(vreg_23_13), .right(vreg_25_13), .up(vreg_24_14), .down(vreg_24_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_13), .sw(sw));
	wire signed[17:0] vwire_24_14;
	reg signed[17:0] vreg_24_14;
	node n24_14(.left(vreg_23_14), .right(vreg_25_14), .up(vreg_24_15), .down(vreg_24_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_14), .sw(sw));
	wire signed[17:0] vwire_24_15;
	reg signed[17:0] vreg_24_15;
	node n24_15(.left(vreg_23_15), .right(vreg_25_15), .up(vreg_24_16), .down(vreg_24_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_15), .sw(sw));
	wire signed[17:0] vwire_24_16;
	reg signed[17:0] vreg_24_16;
	node n24_16(.left(vreg_23_16), .right(vreg_25_16), .up(vreg_24_17), .down(vreg_24_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_16), .sw(sw));
	wire signed[17:0] vwire_24_17;
	reg signed[17:0] vreg_24_17;
	node n24_17(.left(vreg_23_17), .right(vreg_25_17), .up(vreg_24_18), .down(vreg_24_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_17), .sw(sw));
	wire signed[17:0] vwire_24_18;
	reg signed[17:0] vreg_24_18;
	node n24_18(.left(vreg_23_18), .right(vreg_25_18), .up(vreg_24_19), .down(vreg_24_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_18), .sw(sw));
	wire signed[17:0] vwire_24_19;
	reg signed[17:0] vreg_24_19;
	node n24_19(.left(vreg_23_19), .right(vreg_25_19), .up(vreg_24_20), .down(vreg_24_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_19), .sw(sw));
	wire signed[17:0] vwire_24_20;
	reg signed[17:0] vreg_24_20;
	node n24_20(.left(vreg_23_20), .right(vreg_25_20), .up(vreg_24_21), .down(vreg_24_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_20), .sw(sw));
	wire signed[17:0] vwire_24_21;
	reg signed[17:0] vreg_24_21;
	node n24_21(.left(vreg_23_21), .right(vreg_25_21), .up(vreg_24_22), .down(vreg_24_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_21), .sw(sw));
	wire signed[17:0] vwire_24_22;
	reg signed[17:0] vreg_24_22;
	node n24_22(.left(vreg_23_22), .right(vreg_25_22), .up(vreg_24_23), .down(vreg_24_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_22), .sw(sw));
	wire signed[17:0] vwire_24_23;
	reg signed[17:0] vreg_24_23;
	node n24_23(.left(vreg_23_23), .right(vreg_25_23), .up(vreg_24_24), .down(vreg_24_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_23), .sw(sw));
	wire signed[17:0] vwire_24_24;
	reg signed[17:0] vreg_24_24;
	node n24_24(.left(vreg_23_24), .right(vreg_25_24), .up(vreg_24_25), .down(vreg_24_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_24), .sw(sw));
	wire signed[17:0] vwire_24_25;
	reg signed[17:0] vreg_24_25;
	node n24_25(.left(vreg_23_25), .right(vreg_25_25), .up(vreg_24_26), .down(vreg_24_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_25), .sw(sw));
	wire signed[17:0] vwire_24_26;
	reg signed[17:0] vreg_24_26;
	node n24_26(.left(vreg_23_26), .right(vreg_25_26), .up(vreg_24_27), .down(vreg_24_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_26), .sw(sw));
	wire signed[17:0] vwire_24_27;
	reg signed[17:0] vreg_24_27;
	node n24_27(.left(vreg_23_27), .right(vreg_25_27), .up(vreg_24_28), .down(vreg_24_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_27), .sw(sw));
	wire signed[17:0] vwire_24_28;
	reg signed[17:0] vreg_24_28;
	node n24_28(.left(vreg_23_28), .right(vreg_25_28), .up(vreg_24_29), .down(vreg_24_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_28), .sw(sw));
	wire signed[17:0] vwire_24_29;
	reg signed[17:0] vreg_24_29;
	node n24_29(.left(vreg_23_29), .right(vreg_25_29), .up(vreg_24_30), .down(vreg_24_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_29), .sw(sw));
	wire signed[17:0] vwire_24_30;
	reg signed[17:0] vreg_24_30;
	node n24_30(.left(vreg_23_30), .right(vreg_25_30), .up(vreg_24_31), .down(vreg_24_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_30), .sw(sw));
	wire signed[17:0] vwire_24_31;
	reg signed[17:0] vreg_24_31;
	node n24_31(.left(vreg_23_31), .right(vreg_25_31), .up(vreg_24_32), .down(vreg_24_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_31), .sw(sw));
	wire signed[17:0] vwire_24_32;
	reg signed[17:0] vreg_24_32;
	node n24_32(.left(vreg_23_32), .right(vreg_25_32), .up(vreg_24_33), .down(vreg_24_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_32), .sw(sw));
	wire signed[17:0] vwire_24_33;
	reg signed[17:0] vreg_24_33;
	node n24_33(.left(vreg_23_33), .right(vreg_25_33), .up(vreg_24_34), .down(vreg_24_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_33), .sw(sw));
	wire signed[17:0] vwire_24_34;
	reg signed[17:0] vreg_24_34;
	node n24_34(.left(vreg_23_34), .right(vreg_25_34), .up(vreg_24_35), .down(vreg_24_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_34), .sw(sw));
	wire signed[17:0] vwire_24_35;
	reg signed[17:0] vreg_24_35;
	node n24_35(.left(vreg_23_35), .right(vreg_25_35), .up(vreg_24_36), .down(vreg_24_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_35), .sw(sw));
	wire signed[17:0] vwire_24_36;
	reg signed[17:0] vreg_24_36;
	node n24_36(.left(vreg_23_36), .right(vreg_25_36), .up(vreg_24_37), .down(vreg_24_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_36), .sw(sw));
	wire signed[17:0] vwire_24_37;
	reg signed[17:0] vreg_24_37;
	node n24_37(.left(vreg_23_37), .right(vreg_25_37), .up(vreg_24_38), .down(vreg_24_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_37), .sw(sw));
	wire signed[17:0] vwire_24_38;
	reg signed[17:0] vreg_24_38;
	node n24_38(.left(vreg_23_38), .right(vreg_25_38), .up(vreg_24_39), .down(vreg_24_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_38), .sw(sw));
	wire signed[17:0] vwire_24_39;
	reg signed[17:0] vreg_24_39;
	node n24_39(.left(vreg_23_39), .right(vreg_25_39), .up(vreg_24_40), .down(vreg_24_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_39), .sw(sw));
	wire signed[17:0] vwire_24_40;
	reg signed[17:0] vreg_24_40;
	node n24_40(.left(vreg_23_40), .right(vreg_25_40), .up(vreg_24_41), .down(vreg_24_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_40), .sw(sw));
	wire signed[17:0] vwire_24_41;
	reg signed[17:0] vreg_24_41;
	node n24_41(.left(vreg_23_41), .right(vreg_25_41), .up(vreg_24_42), .down(vreg_24_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_41), .sw(sw));
	wire signed[17:0] vwire_24_42;
	reg signed[17:0] vreg_24_42;
	node n24_42(.left(vreg_23_42), .right(vreg_25_42), .up(vreg_24_43), .down(vreg_24_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_42), .sw(sw));
	wire signed[17:0] vwire_24_43;
	reg signed[17:0] vreg_24_43;
	node n24_43(.left(vreg_23_43), .right(vreg_25_43), .up(vreg_24_44), .down(vreg_24_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_43), .sw(sw));
	wire signed[17:0] vwire_24_44;
	reg signed[17:0] vreg_24_44;
	node n24_44(.left(vreg_23_44), .right(vreg_25_44), .up(vreg_24_45), .down(vreg_24_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_44), .sw(sw));
	wire signed[17:0] vwire_24_45;
	reg signed[17:0] vreg_24_45;
	node n24_45(.left(vreg_23_45), .right(vreg_25_45), .up(vreg_24_46), .down(vreg_24_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_45), .sw(sw));
	wire signed[17:0] vwire_24_46;
	reg signed[17:0] vreg_24_46;
	node n24_46(.left(vreg_23_46), .right(vreg_25_46), .up(vreg_24_47), .down(vreg_24_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_46), .sw(sw));
	wire signed[17:0] vwire_24_47;
	reg signed[17:0] vreg_24_47;
	node n24_47(.left(vreg_23_47), .right(vreg_25_47), .up(vreg_24_48), .down(vreg_24_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_47), .sw(sw));
	wire signed[17:0] vwire_24_48;
	reg signed[17:0] vreg_24_48;
	node n24_48(.left(vreg_23_48), .right(vreg_25_48), .up(vreg_24_49), .down(vreg_24_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_48), .sw(sw));
	wire signed[17:0] vwire_24_49;
	reg signed[17:0] vreg_24_49;
	node n24_49(.left(vreg_23_49), .right(vreg_25_49), .up(18'b0), .down(vreg_24_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_24_49), .sw(sw));
	wire signed[17:0] vwire_25_0;
	reg signed[17:0] vreg_25_0;
	node n25_0(.left(vreg_24_0), .right(vreg_26_0), .up(vreg_25_1), .down(vreg_25_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_0), .sw(sw));
	wire signed[17:0] vwire_25_1;
	reg signed[17:0] vreg_25_1;
	node n25_1(.left(vreg_24_1), .right(vreg_26_1), .up(vreg_25_2), .down(vreg_25_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_1), .sw(sw));
	wire signed[17:0] vwire_25_2;
	reg signed[17:0] vreg_25_2;
	node n25_2(.left(vreg_24_2), .right(vreg_26_2), .up(vreg_25_3), .down(vreg_25_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_2), .sw(sw));
	wire signed[17:0] vwire_25_3;
	reg signed[17:0] vreg_25_3;
	node n25_3(.left(vreg_24_3), .right(vreg_26_3), .up(vreg_25_4), .down(vreg_25_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_3), .sw(sw));
	wire signed[17:0] vwire_25_4;
	reg signed[17:0] vreg_25_4;
	node n25_4(.left(vreg_24_4), .right(vreg_26_4), .up(vreg_25_5), .down(vreg_25_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_4), .sw(sw));
	wire signed[17:0] vwire_25_5;
	reg signed[17:0] vreg_25_5;
	node n25_5(.left(vreg_24_5), .right(vreg_26_5), .up(vreg_25_6), .down(vreg_25_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_5), .sw(sw));
	wire signed[17:0] vwire_25_6;
	reg signed[17:0] vreg_25_6;
	node n25_6(.left(vreg_24_6), .right(vreg_26_6), .up(vreg_25_7), .down(vreg_25_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_6), .sw(sw));
	wire signed[17:0] vwire_25_7;
	reg signed[17:0] vreg_25_7;
	node n25_7(.left(vreg_24_7), .right(vreg_26_7), .up(vreg_25_8), .down(vreg_25_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_7), .sw(sw));
	wire signed[17:0] vwire_25_8;
	reg signed[17:0] vreg_25_8;
	node n25_8(.left(vreg_24_8), .right(vreg_26_8), .up(vreg_25_9), .down(vreg_25_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_8), .sw(sw));
	wire signed[17:0] vwire_25_9;
	reg signed[17:0] vreg_25_9;
	node n25_9(.left(vreg_24_9), .right(vreg_26_9), .up(vreg_25_10), .down(vreg_25_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_9), .sw(sw));
	wire signed[17:0] vwire_25_10;
	reg signed[17:0] vreg_25_10;
	node n25_10(.left(vreg_24_10), .right(vreg_26_10), .up(vreg_25_11), .down(vreg_25_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_10), .sw(sw));
	wire signed[17:0] vwire_25_11;
	reg signed[17:0] vreg_25_11;
	node n25_11(.left(vreg_24_11), .right(vreg_26_11), .up(vreg_25_12), .down(vreg_25_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_11), .sw(sw));
	wire signed[17:0] vwire_25_12;
	reg signed[17:0] vreg_25_12;
	node n25_12(.left(vreg_24_12), .right(vreg_26_12), .up(vreg_25_13), .down(vreg_25_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_12), .sw(sw));
	wire signed[17:0] vwire_25_13;
	reg signed[17:0] vreg_25_13;
	node n25_13(.left(vreg_24_13), .right(vreg_26_13), .up(vreg_25_14), .down(vreg_25_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_13), .sw(sw));
	wire signed[17:0] vwire_25_14;
	reg signed[17:0] vreg_25_14;
	node n25_14(.left(vreg_24_14), .right(vreg_26_14), .up(vreg_25_15), .down(vreg_25_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_14), .sw(sw));
	wire signed[17:0] vwire_25_15;
	reg signed[17:0] vreg_25_15;
	node n25_15(.left(vreg_24_15), .right(vreg_26_15), .up(vreg_25_16), .down(vreg_25_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_15), .sw(sw));
	wire signed[17:0] vwire_25_16;
	reg signed[17:0] vreg_25_16;
	node n25_16(.left(vreg_24_16), .right(vreg_26_16), .up(vreg_25_17), .down(vreg_25_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_16), .sw(sw));
	wire signed[17:0] vwire_25_17;
	reg signed[17:0] vreg_25_17;
	node n25_17(.left(vreg_24_17), .right(vreg_26_17), .up(vreg_25_18), .down(vreg_25_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_17), .sw(sw));
	wire signed[17:0] vwire_25_18;
	reg signed[17:0] vreg_25_18;
	node n25_18(.left(vreg_24_18), .right(vreg_26_18), .up(vreg_25_19), .down(vreg_25_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_18), .sw(sw));
	wire signed[17:0] vwire_25_19;
	reg signed[17:0] vreg_25_19;
	node n25_19(.left(vreg_24_19), .right(vreg_26_19), .up(vreg_25_20), .down(vreg_25_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_19), .sw(sw));
	wire signed[17:0] vwire_25_20;
	reg signed[17:0] vreg_25_20;
	node n25_20(.left(vreg_24_20), .right(vreg_26_20), .up(vreg_25_21), .down(vreg_25_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_20), .sw(sw));
	wire signed[17:0] vwire_25_21;
	reg signed[17:0] vreg_25_21;
	node n25_21(.left(vreg_24_21), .right(vreg_26_21), .up(vreg_25_22), .down(vreg_25_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_21), .sw(sw));
	wire signed[17:0] vwire_25_22;
	reg signed[17:0] vreg_25_22;
	node n25_22(.left(vreg_24_22), .right(vreg_26_22), .up(vreg_25_23), .down(vreg_25_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_22), .sw(sw));
	wire signed[17:0] vwire_25_23;
	reg signed[17:0] vreg_25_23;
	node n25_23(.left(vreg_24_23), .right(vreg_26_23), .up(vreg_25_24), .down(vreg_25_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_23), .sw(sw));
	wire signed[17:0] vwire_25_24;
	reg signed[17:0] vreg_25_24;
	node n25_24(.left(vreg_24_24), .right(vreg_26_24), .up(vreg_25_25), .down(vreg_25_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_24), .sw(sw));
	wire signed[17:0] vwire_25_25;
	reg signed[17:0] vreg_25_25;
	node n25_25(.left(vreg_24_25), .right(vreg_26_25), .up(vreg_25_26), .down(vreg_25_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_25), .sw(sw));
	wire signed[17:0] vwire_25_26;
	reg signed[17:0] vreg_25_26;
	node n25_26(.left(vreg_24_26), .right(vreg_26_26), .up(vreg_25_27), .down(vreg_25_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_26), .sw(sw));
	wire signed[17:0] vwire_25_27;
	reg signed[17:0] vreg_25_27;
	node n25_27(.left(vreg_24_27), .right(vreg_26_27), .up(vreg_25_28), .down(vreg_25_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_27), .sw(sw));
	wire signed[17:0] vwire_25_28;
	reg signed[17:0] vreg_25_28;
	node n25_28(.left(vreg_24_28), .right(vreg_26_28), .up(vreg_25_29), .down(vreg_25_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_28), .sw(sw));
	wire signed[17:0] vwire_25_29;
	reg signed[17:0] vreg_25_29;
	node n25_29(.left(vreg_24_29), .right(vreg_26_29), .up(vreg_25_30), .down(vreg_25_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_29), .sw(sw));
	wire signed[17:0] vwire_25_30;
	reg signed[17:0] vreg_25_30;
	node n25_30(.left(vreg_24_30), .right(vreg_26_30), .up(vreg_25_31), .down(vreg_25_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_30), .sw(sw));
	wire signed[17:0] vwire_25_31;
	reg signed[17:0] vreg_25_31;
	node n25_31(.left(vreg_24_31), .right(vreg_26_31), .up(vreg_25_32), .down(vreg_25_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_31), .sw(sw));
	wire signed[17:0] vwire_25_32;
	reg signed[17:0] vreg_25_32;
	node n25_32(.left(vreg_24_32), .right(vreg_26_32), .up(vreg_25_33), .down(vreg_25_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_32), .sw(sw));
	wire signed[17:0] vwire_25_33;
	reg signed[17:0] vreg_25_33;
	node n25_33(.left(vreg_24_33), .right(vreg_26_33), .up(vreg_25_34), .down(vreg_25_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_33), .sw(sw));
	wire signed[17:0] vwire_25_34;
	reg signed[17:0] vreg_25_34;
	node n25_34(.left(vreg_24_34), .right(vreg_26_34), .up(vreg_25_35), .down(vreg_25_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_34), .sw(sw));
	wire signed[17:0] vwire_25_35;
	reg signed[17:0] vreg_25_35;
	node n25_35(.left(vreg_24_35), .right(vreg_26_35), .up(vreg_25_36), .down(vreg_25_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_35), .sw(sw));
	wire signed[17:0] vwire_25_36;
	reg signed[17:0] vreg_25_36;
	node n25_36(.left(vreg_24_36), .right(vreg_26_36), .up(vreg_25_37), .down(vreg_25_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_36), .sw(sw));
	wire signed[17:0] vwire_25_37;
	reg signed[17:0] vreg_25_37;
	node n25_37(.left(vreg_24_37), .right(vreg_26_37), .up(vreg_25_38), .down(vreg_25_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_37), .sw(sw));
	wire signed[17:0] vwire_25_38;
	reg signed[17:0] vreg_25_38;
	node n25_38(.left(vreg_24_38), .right(vreg_26_38), .up(vreg_25_39), .down(vreg_25_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_38), .sw(sw));
	wire signed[17:0] vwire_25_39;
	reg signed[17:0] vreg_25_39;
	node n25_39(.left(vreg_24_39), .right(vreg_26_39), .up(vreg_25_40), .down(vreg_25_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_39), .sw(sw));
	wire signed[17:0] vwire_25_40;
	reg signed[17:0] vreg_25_40;
	node n25_40(.left(vreg_24_40), .right(vreg_26_40), .up(vreg_25_41), .down(vreg_25_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_40), .sw(sw));
	wire signed[17:0] vwire_25_41;
	reg signed[17:0] vreg_25_41;
	node n25_41(.left(vreg_24_41), .right(vreg_26_41), .up(vreg_25_42), .down(vreg_25_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_41), .sw(sw));
	wire signed[17:0] vwire_25_42;
	reg signed[17:0] vreg_25_42;
	node n25_42(.left(vreg_24_42), .right(vreg_26_42), .up(vreg_25_43), .down(vreg_25_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_42), .sw(sw));
	wire signed[17:0] vwire_25_43;
	reg signed[17:0] vreg_25_43;
	node n25_43(.left(vreg_24_43), .right(vreg_26_43), .up(vreg_25_44), .down(vreg_25_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_43), .sw(sw));
	wire signed[17:0] vwire_25_44;
	reg signed[17:0] vreg_25_44;
	node n25_44(.left(vreg_24_44), .right(vreg_26_44), .up(vreg_25_45), .down(vreg_25_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_44), .sw(sw));
	wire signed[17:0] vwire_25_45;
	reg signed[17:0] vreg_25_45;
	node n25_45(.left(vreg_24_45), .right(vreg_26_45), .up(vreg_25_46), .down(vreg_25_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_45), .sw(sw));
	wire signed[17:0] vwire_25_46;
	reg signed[17:0] vreg_25_46;
	node n25_46(.left(vreg_24_46), .right(vreg_26_46), .up(vreg_25_47), .down(vreg_25_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_46), .sw(sw));
	wire signed[17:0] vwire_25_47;
	reg signed[17:0] vreg_25_47;
	node n25_47(.left(vreg_24_47), .right(vreg_26_47), .up(vreg_25_48), .down(vreg_25_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_47), .sw(sw));
	wire signed[17:0] vwire_25_48;
	reg signed[17:0] vreg_25_48;
	node n25_48(.left(vreg_24_48), .right(vreg_26_48), .up(vreg_25_49), .down(vreg_25_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_48), .sw(sw));
	wire signed[17:0] vwire_25_49;
	reg signed[17:0] vreg_25_49;
	node n25_49(.left(vreg_24_49), .right(vreg_26_49), .up(18'b0), .down(vreg_25_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_25_49), .sw(sw));
	wire signed[17:0] vwire_26_0;
	reg signed[17:0] vreg_26_0;
	node n26_0(.left(vreg_25_0), .right(vreg_27_0), .up(vreg_26_1), .down(vreg_26_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_0), .sw(sw));
	wire signed[17:0] vwire_26_1;
	reg signed[17:0] vreg_26_1;
	node n26_1(.left(vreg_25_1), .right(vreg_27_1), .up(vreg_26_2), .down(vreg_26_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_1), .sw(sw));
	wire signed[17:0] vwire_26_2;
	reg signed[17:0] vreg_26_2;
	node n26_2(.left(vreg_25_2), .right(vreg_27_2), .up(vreg_26_3), .down(vreg_26_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_2), .sw(sw));
	wire signed[17:0] vwire_26_3;
	reg signed[17:0] vreg_26_3;
	node n26_3(.left(vreg_25_3), .right(vreg_27_3), .up(vreg_26_4), .down(vreg_26_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_3), .sw(sw));
	wire signed[17:0] vwire_26_4;
	reg signed[17:0] vreg_26_4;
	node n26_4(.left(vreg_25_4), .right(vreg_27_4), .up(vreg_26_5), .down(vreg_26_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_4), .sw(sw));
	wire signed[17:0] vwire_26_5;
	reg signed[17:0] vreg_26_5;
	node n26_5(.left(vreg_25_5), .right(vreg_27_5), .up(vreg_26_6), .down(vreg_26_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_5), .sw(sw));
	wire signed[17:0] vwire_26_6;
	reg signed[17:0] vreg_26_6;
	node n26_6(.left(vreg_25_6), .right(vreg_27_6), .up(vreg_26_7), .down(vreg_26_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_6), .sw(sw));
	wire signed[17:0] vwire_26_7;
	reg signed[17:0] vreg_26_7;
	node n26_7(.left(vreg_25_7), .right(vreg_27_7), .up(vreg_26_8), .down(vreg_26_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_7), .sw(sw));
	wire signed[17:0] vwire_26_8;
	reg signed[17:0] vreg_26_8;
	node n26_8(.left(vreg_25_8), .right(vreg_27_8), .up(vreg_26_9), .down(vreg_26_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_8), .sw(sw));
	wire signed[17:0] vwire_26_9;
	reg signed[17:0] vreg_26_9;
	node n26_9(.left(vreg_25_9), .right(vreg_27_9), .up(vreg_26_10), .down(vreg_26_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_9), .sw(sw));
	wire signed[17:0] vwire_26_10;
	reg signed[17:0] vreg_26_10;
	node n26_10(.left(vreg_25_10), .right(vreg_27_10), .up(vreg_26_11), .down(vreg_26_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_10), .sw(sw));
	wire signed[17:0] vwire_26_11;
	reg signed[17:0] vreg_26_11;
	node n26_11(.left(vreg_25_11), .right(vreg_27_11), .up(vreg_26_12), .down(vreg_26_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_11), .sw(sw));
	wire signed[17:0] vwire_26_12;
	reg signed[17:0] vreg_26_12;
	node n26_12(.left(vreg_25_12), .right(vreg_27_12), .up(vreg_26_13), .down(vreg_26_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_12), .sw(sw));
	wire signed[17:0] vwire_26_13;
	reg signed[17:0] vreg_26_13;
	node n26_13(.left(vreg_25_13), .right(vreg_27_13), .up(vreg_26_14), .down(vreg_26_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_13), .sw(sw));
	wire signed[17:0] vwire_26_14;
	reg signed[17:0] vreg_26_14;
	node n26_14(.left(vreg_25_14), .right(vreg_27_14), .up(vreg_26_15), .down(vreg_26_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_14), .sw(sw));
	wire signed[17:0] vwire_26_15;
	reg signed[17:0] vreg_26_15;
	node n26_15(.left(vreg_25_15), .right(vreg_27_15), .up(vreg_26_16), .down(vreg_26_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_15), .sw(sw));
	wire signed[17:0] vwire_26_16;
	reg signed[17:0] vreg_26_16;
	node n26_16(.left(vreg_25_16), .right(vreg_27_16), .up(vreg_26_17), .down(vreg_26_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_16), .sw(sw));
	wire signed[17:0] vwire_26_17;
	reg signed[17:0] vreg_26_17;
	node n26_17(.left(vreg_25_17), .right(vreg_27_17), .up(vreg_26_18), .down(vreg_26_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_17), .sw(sw));
	wire signed[17:0] vwire_26_18;
	reg signed[17:0] vreg_26_18;
	node n26_18(.left(vreg_25_18), .right(vreg_27_18), .up(vreg_26_19), .down(vreg_26_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_18), .sw(sw));
	wire signed[17:0] vwire_26_19;
	reg signed[17:0] vreg_26_19;
	node n26_19(.left(vreg_25_19), .right(vreg_27_19), .up(vreg_26_20), .down(vreg_26_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_19), .sw(sw));
	wire signed[17:0] vwire_26_20;
	reg signed[17:0] vreg_26_20;
	node n26_20(.left(vreg_25_20), .right(vreg_27_20), .up(vreg_26_21), .down(vreg_26_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_20), .sw(sw));
	wire signed[17:0] vwire_26_21;
	reg signed[17:0] vreg_26_21;
	node n26_21(.left(vreg_25_21), .right(vreg_27_21), .up(vreg_26_22), .down(vreg_26_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_21), .sw(sw));
	wire signed[17:0] vwire_26_22;
	reg signed[17:0] vreg_26_22;
	node n26_22(.left(vreg_25_22), .right(vreg_27_22), .up(vreg_26_23), .down(vreg_26_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_22), .sw(sw));
	wire signed[17:0] vwire_26_23;
	reg signed[17:0] vreg_26_23;
	node n26_23(.left(vreg_25_23), .right(vreg_27_23), .up(vreg_26_24), .down(vreg_26_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_23), .sw(sw));
	wire signed[17:0] vwire_26_24;
	reg signed[17:0] vreg_26_24;
	node n26_24(.left(vreg_25_24), .right(vreg_27_24), .up(vreg_26_25), .down(vreg_26_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_24), .sw(sw));
	wire signed[17:0] vwire_26_25;
	reg signed[17:0] vreg_26_25;
	node n26_25(.left(vreg_25_25), .right(vreg_27_25), .up(vreg_26_26), .down(vreg_26_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_25), .sw(sw));
	wire signed[17:0] vwire_26_26;
	reg signed[17:0] vreg_26_26;
	node n26_26(.left(vreg_25_26), .right(vreg_27_26), .up(vreg_26_27), .down(vreg_26_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_26), .sw(sw));
	wire signed[17:0] vwire_26_27;
	reg signed[17:0] vreg_26_27;
	node n26_27(.left(vreg_25_27), .right(vreg_27_27), .up(vreg_26_28), .down(vreg_26_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_27), .sw(sw));
	wire signed[17:0] vwire_26_28;
	reg signed[17:0] vreg_26_28;
	node n26_28(.left(vreg_25_28), .right(vreg_27_28), .up(vreg_26_29), .down(vreg_26_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_28), .sw(sw));
	wire signed[17:0] vwire_26_29;
	reg signed[17:0] vreg_26_29;
	node n26_29(.left(vreg_25_29), .right(vreg_27_29), .up(vreg_26_30), .down(vreg_26_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_29), .sw(sw));
	wire signed[17:0] vwire_26_30;
	reg signed[17:0] vreg_26_30;
	node n26_30(.left(vreg_25_30), .right(vreg_27_30), .up(vreg_26_31), .down(vreg_26_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_30), .sw(sw));
	wire signed[17:0] vwire_26_31;
	reg signed[17:0] vreg_26_31;
	node n26_31(.left(vreg_25_31), .right(vreg_27_31), .up(vreg_26_32), .down(vreg_26_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_31), .sw(sw));
	wire signed[17:0] vwire_26_32;
	reg signed[17:0] vreg_26_32;
	node n26_32(.left(vreg_25_32), .right(vreg_27_32), .up(vreg_26_33), .down(vreg_26_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_32), .sw(sw));
	wire signed[17:0] vwire_26_33;
	reg signed[17:0] vreg_26_33;
	node n26_33(.left(vreg_25_33), .right(vreg_27_33), .up(vreg_26_34), .down(vreg_26_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_33), .sw(sw));
	wire signed[17:0] vwire_26_34;
	reg signed[17:0] vreg_26_34;
	node n26_34(.left(vreg_25_34), .right(vreg_27_34), .up(vreg_26_35), .down(vreg_26_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_34), .sw(sw));
	wire signed[17:0] vwire_26_35;
	reg signed[17:0] vreg_26_35;
	node n26_35(.left(vreg_25_35), .right(vreg_27_35), .up(vreg_26_36), .down(vreg_26_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_35), .sw(sw));
	wire signed[17:0] vwire_26_36;
	reg signed[17:0] vreg_26_36;
	node n26_36(.left(vreg_25_36), .right(vreg_27_36), .up(vreg_26_37), .down(vreg_26_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_36), .sw(sw));
	wire signed[17:0] vwire_26_37;
	reg signed[17:0] vreg_26_37;
	node n26_37(.left(vreg_25_37), .right(vreg_27_37), .up(vreg_26_38), .down(vreg_26_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_37), .sw(sw));
	wire signed[17:0] vwire_26_38;
	reg signed[17:0] vreg_26_38;
	node n26_38(.left(vreg_25_38), .right(vreg_27_38), .up(vreg_26_39), .down(vreg_26_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_38), .sw(sw));
	wire signed[17:0] vwire_26_39;
	reg signed[17:0] vreg_26_39;
	node n26_39(.left(vreg_25_39), .right(vreg_27_39), .up(vreg_26_40), .down(vreg_26_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_39), .sw(sw));
	wire signed[17:0] vwire_26_40;
	reg signed[17:0] vreg_26_40;
	node n26_40(.left(vreg_25_40), .right(vreg_27_40), .up(vreg_26_41), .down(vreg_26_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_40), .sw(sw));
	wire signed[17:0] vwire_26_41;
	reg signed[17:0] vreg_26_41;
	node n26_41(.left(vreg_25_41), .right(vreg_27_41), .up(vreg_26_42), .down(vreg_26_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_41), .sw(sw));
	wire signed[17:0] vwire_26_42;
	reg signed[17:0] vreg_26_42;
	node n26_42(.left(vreg_25_42), .right(vreg_27_42), .up(vreg_26_43), .down(vreg_26_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_42), .sw(sw));
	wire signed[17:0] vwire_26_43;
	reg signed[17:0] vreg_26_43;
	node n26_43(.left(vreg_25_43), .right(vreg_27_43), .up(vreg_26_44), .down(vreg_26_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_43), .sw(sw));
	wire signed[17:0] vwire_26_44;
	reg signed[17:0] vreg_26_44;
	node n26_44(.left(vreg_25_44), .right(vreg_27_44), .up(vreg_26_45), .down(vreg_26_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_44), .sw(sw));
	wire signed[17:0] vwire_26_45;
	reg signed[17:0] vreg_26_45;
	node n26_45(.left(vreg_25_45), .right(vreg_27_45), .up(vreg_26_46), .down(vreg_26_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_45), .sw(sw));
	wire signed[17:0] vwire_26_46;
	reg signed[17:0] vreg_26_46;
	node n26_46(.left(vreg_25_46), .right(vreg_27_46), .up(vreg_26_47), .down(vreg_26_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_46), .sw(sw));
	wire signed[17:0] vwire_26_47;
	reg signed[17:0] vreg_26_47;
	node n26_47(.left(vreg_25_47), .right(vreg_27_47), .up(vreg_26_48), .down(vreg_26_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_47), .sw(sw));
	wire signed[17:0] vwire_26_48;
	reg signed[17:0] vreg_26_48;
	node n26_48(.left(vreg_25_48), .right(vreg_27_48), .up(vreg_26_49), .down(vreg_26_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_48), .sw(sw));
	wire signed[17:0] vwire_26_49;
	reg signed[17:0] vreg_26_49;
	node n26_49(.left(vreg_25_49), .right(vreg_27_49), .up(18'b0), .down(vreg_26_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_26_49), .sw(sw));
	wire signed[17:0] vwire_27_0;
	reg signed[17:0] vreg_27_0;
	node n27_0(.left(vreg_26_0), .right(vreg_28_0), .up(vreg_27_1), .down(vreg_27_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_0), .sw(sw));
	wire signed[17:0] vwire_27_1;
	reg signed[17:0] vreg_27_1;
	node n27_1(.left(vreg_26_1), .right(vreg_28_1), .up(vreg_27_2), .down(vreg_27_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_1), .sw(sw));
	wire signed[17:0] vwire_27_2;
	reg signed[17:0] vreg_27_2;
	node n27_2(.left(vreg_26_2), .right(vreg_28_2), .up(vreg_27_3), .down(vreg_27_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_2), .sw(sw));
	wire signed[17:0] vwire_27_3;
	reg signed[17:0] vreg_27_3;
	node n27_3(.left(vreg_26_3), .right(vreg_28_3), .up(vreg_27_4), .down(vreg_27_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_3), .sw(sw));
	wire signed[17:0] vwire_27_4;
	reg signed[17:0] vreg_27_4;
	node n27_4(.left(vreg_26_4), .right(vreg_28_4), .up(vreg_27_5), .down(vreg_27_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_4), .sw(sw));
	wire signed[17:0] vwire_27_5;
	reg signed[17:0] vreg_27_5;
	node n27_5(.left(vreg_26_5), .right(vreg_28_5), .up(vreg_27_6), .down(vreg_27_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_5), .sw(sw));
	wire signed[17:0] vwire_27_6;
	reg signed[17:0] vreg_27_6;
	node n27_6(.left(vreg_26_6), .right(vreg_28_6), .up(vreg_27_7), .down(vreg_27_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_6), .sw(sw));
	wire signed[17:0] vwire_27_7;
	reg signed[17:0] vreg_27_7;
	node n27_7(.left(vreg_26_7), .right(vreg_28_7), .up(vreg_27_8), .down(vreg_27_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_7), .sw(sw));
	wire signed[17:0] vwire_27_8;
	reg signed[17:0] vreg_27_8;
	node n27_8(.left(vreg_26_8), .right(vreg_28_8), .up(vreg_27_9), .down(vreg_27_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_8), .sw(sw));
	wire signed[17:0] vwire_27_9;
	reg signed[17:0] vreg_27_9;
	node n27_9(.left(vreg_26_9), .right(vreg_28_9), .up(vreg_27_10), .down(vreg_27_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_9), .sw(sw));
	wire signed[17:0] vwire_27_10;
	reg signed[17:0] vreg_27_10;
	node n27_10(.left(vreg_26_10), .right(vreg_28_10), .up(vreg_27_11), .down(vreg_27_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_10), .sw(sw));
	wire signed[17:0] vwire_27_11;
	reg signed[17:0] vreg_27_11;
	node n27_11(.left(vreg_26_11), .right(vreg_28_11), .up(vreg_27_12), .down(vreg_27_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_11), .sw(sw));
	wire signed[17:0] vwire_27_12;
	reg signed[17:0] vreg_27_12;
	node n27_12(.left(vreg_26_12), .right(vreg_28_12), .up(vreg_27_13), .down(vreg_27_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_12), .sw(sw));
	wire signed[17:0] vwire_27_13;
	reg signed[17:0] vreg_27_13;
	node n27_13(.left(vreg_26_13), .right(vreg_28_13), .up(vreg_27_14), .down(vreg_27_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_13), .sw(sw));
	wire signed[17:0] vwire_27_14;
	reg signed[17:0] vreg_27_14;
	node n27_14(.left(vreg_26_14), .right(vreg_28_14), .up(vreg_27_15), .down(vreg_27_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_14), .sw(sw));
	wire signed[17:0] vwire_27_15;
	reg signed[17:0] vreg_27_15;
	node n27_15(.left(vreg_26_15), .right(vreg_28_15), .up(vreg_27_16), .down(vreg_27_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_15), .sw(sw));
	wire signed[17:0] vwire_27_16;
	reg signed[17:0] vreg_27_16;
	node n27_16(.left(vreg_26_16), .right(vreg_28_16), .up(vreg_27_17), .down(vreg_27_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_16), .sw(sw));
	wire signed[17:0] vwire_27_17;
	reg signed[17:0] vreg_27_17;
	node n27_17(.left(vreg_26_17), .right(vreg_28_17), .up(vreg_27_18), .down(vreg_27_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_17), .sw(sw));
	wire signed[17:0] vwire_27_18;
	reg signed[17:0] vreg_27_18;
	node n27_18(.left(vreg_26_18), .right(vreg_28_18), .up(vreg_27_19), .down(vreg_27_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_18), .sw(sw));
	wire signed[17:0] vwire_27_19;
	reg signed[17:0] vreg_27_19;
	node n27_19(.left(vreg_26_19), .right(vreg_28_19), .up(vreg_27_20), .down(vreg_27_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_19), .sw(sw));
	wire signed[17:0] vwire_27_20;
	reg signed[17:0] vreg_27_20;
	node n27_20(.left(vreg_26_20), .right(vreg_28_20), .up(vreg_27_21), .down(vreg_27_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_20), .sw(sw));
	wire signed[17:0] vwire_27_21;
	reg signed[17:0] vreg_27_21;
	node n27_21(.left(vreg_26_21), .right(vreg_28_21), .up(vreg_27_22), .down(vreg_27_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_21), .sw(sw));
	wire signed[17:0] vwire_27_22;
	reg signed[17:0] vreg_27_22;
	node n27_22(.left(vreg_26_22), .right(vreg_28_22), .up(vreg_27_23), .down(vreg_27_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_22), .sw(sw));
	wire signed[17:0] vwire_27_23;
	reg signed[17:0] vreg_27_23;
	node n27_23(.left(vreg_26_23), .right(vreg_28_23), .up(vreg_27_24), .down(vreg_27_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_23), .sw(sw));
	wire signed[17:0] vwire_27_24;
	reg signed[17:0] vreg_27_24;
	node n27_24(.left(vreg_26_24), .right(vreg_28_24), .up(vreg_27_25), .down(vreg_27_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_24), .sw(sw));
	wire signed[17:0] vwire_27_25;
	reg signed[17:0] vreg_27_25;
	node n27_25(.left(vreg_26_25), .right(vreg_28_25), .up(vreg_27_26), .down(vreg_27_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_25), .sw(sw));
	wire signed[17:0] vwire_27_26;
	reg signed[17:0] vreg_27_26;
	node n27_26(.left(vreg_26_26), .right(vreg_28_26), .up(vreg_27_27), .down(vreg_27_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_26), .sw(sw));
	wire signed[17:0] vwire_27_27;
	reg signed[17:0] vreg_27_27;
	node n27_27(.left(vreg_26_27), .right(vreg_28_27), .up(vreg_27_28), .down(vreg_27_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_27), .sw(sw));
	wire signed[17:0] vwire_27_28;
	reg signed[17:0] vreg_27_28;
	node n27_28(.left(vreg_26_28), .right(vreg_28_28), .up(vreg_27_29), .down(vreg_27_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_28), .sw(sw));
	wire signed[17:0] vwire_27_29;
	reg signed[17:0] vreg_27_29;
	node n27_29(.left(vreg_26_29), .right(vreg_28_29), .up(vreg_27_30), .down(vreg_27_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_29), .sw(sw));
	wire signed[17:0] vwire_27_30;
	reg signed[17:0] vreg_27_30;
	node n27_30(.left(vreg_26_30), .right(vreg_28_30), .up(vreg_27_31), .down(vreg_27_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_30), .sw(sw));
	wire signed[17:0] vwire_27_31;
	reg signed[17:0] vreg_27_31;
	node n27_31(.left(vreg_26_31), .right(vreg_28_31), .up(vreg_27_32), .down(vreg_27_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_31), .sw(sw));
	wire signed[17:0] vwire_27_32;
	reg signed[17:0] vreg_27_32;
	node n27_32(.left(vreg_26_32), .right(vreg_28_32), .up(vreg_27_33), .down(vreg_27_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_32), .sw(sw));
	wire signed[17:0] vwire_27_33;
	reg signed[17:0] vreg_27_33;
	node n27_33(.left(vreg_26_33), .right(vreg_28_33), .up(vreg_27_34), .down(vreg_27_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_33), .sw(sw));
	wire signed[17:0] vwire_27_34;
	reg signed[17:0] vreg_27_34;
	node n27_34(.left(vreg_26_34), .right(vreg_28_34), .up(vreg_27_35), .down(vreg_27_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_34), .sw(sw));
	wire signed[17:0] vwire_27_35;
	reg signed[17:0] vreg_27_35;
	node n27_35(.left(vreg_26_35), .right(vreg_28_35), .up(vreg_27_36), .down(vreg_27_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_35), .sw(sw));
	wire signed[17:0] vwire_27_36;
	reg signed[17:0] vreg_27_36;
	node n27_36(.left(vreg_26_36), .right(vreg_28_36), .up(vreg_27_37), .down(vreg_27_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_36), .sw(sw));
	wire signed[17:0] vwire_27_37;
	reg signed[17:0] vreg_27_37;
	node n27_37(.left(vreg_26_37), .right(vreg_28_37), .up(vreg_27_38), .down(vreg_27_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_37), .sw(sw));
	wire signed[17:0] vwire_27_38;
	reg signed[17:0] vreg_27_38;
	node n27_38(.left(vreg_26_38), .right(vreg_28_38), .up(vreg_27_39), .down(vreg_27_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_38), .sw(sw));
	wire signed[17:0] vwire_27_39;
	reg signed[17:0] vreg_27_39;
	node n27_39(.left(vreg_26_39), .right(vreg_28_39), .up(vreg_27_40), .down(vreg_27_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_39), .sw(sw));
	wire signed[17:0] vwire_27_40;
	reg signed[17:0] vreg_27_40;
	node n27_40(.left(vreg_26_40), .right(vreg_28_40), .up(vreg_27_41), .down(vreg_27_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_40), .sw(sw));
	wire signed[17:0] vwire_27_41;
	reg signed[17:0] vreg_27_41;
	node n27_41(.left(vreg_26_41), .right(vreg_28_41), .up(vreg_27_42), .down(vreg_27_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_41), .sw(sw));
	wire signed[17:0] vwire_27_42;
	reg signed[17:0] vreg_27_42;
	node n27_42(.left(vreg_26_42), .right(vreg_28_42), .up(vreg_27_43), .down(vreg_27_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_42), .sw(sw));
	wire signed[17:0] vwire_27_43;
	reg signed[17:0] vreg_27_43;
	node n27_43(.left(vreg_26_43), .right(vreg_28_43), .up(vreg_27_44), .down(vreg_27_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_43), .sw(sw));
	wire signed[17:0] vwire_27_44;
	reg signed[17:0] vreg_27_44;
	node n27_44(.left(vreg_26_44), .right(vreg_28_44), .up(vreg_27_45), .down(vreg_27_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_44), .sw(sw));
	wire signed[17:0] vwire_27_45;
	reg signed[17:0] vreg_27_45;
	node n27_45(.left(vreg_26_45), .right(vreg_28_45), .up(vreg_27_46), .down(vreg_27_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_45), .sw(sw));
	wire signed[17:0] vwire_27_46;
	reg signed[17:0] vreg_27_46;
	node n27_46(.left(vreg_26_46), .right(vreg_28_46), .up(vreg_27_47), .down(vreg_27_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_46), .sw(sw));
	wire signed[17:0] vwire_27_47;
	reg signed[17:0] vreg_27_47;
	node n27_47(.left(vreg_26_47), .right(vreg_28_47), .up(vreg_27_48), .down(vreg_27_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_47), .sw(sw));
	wire signed[17:0] vwire_27_48;
	reg signed[17:0] vreg_27_48;
	node n27_48(.left(vreg_26_48), .right(vreg_28_48), .up(vreg_27_49), .down(vreg_27_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_48), .sw(sw));
	wire signed[17:0] vwire_27_49;
	reg signed[17:0] vreg_27_49;
	node n27_49(.left(vreg_26_49), .right(vreg_28_49), .up(18'b0), .down(vreg_27_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_27_49), .sw(sw));
	wire signed[17:0] vwire_28_0;
	reg signed[17:0] vreg_28_0;
	node n28_0(.left(vreg_27_0), .right(vreg_29_0), .up(vreg_28_1), .down(vreg_28_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_0), .sw(sw));
	wire signed[17:0] vwire_28_1;
	reg signed[17:0] vreg_28_1;
	node n28_1(.left(vreg_27_1), .right(vreg_29_1), .up(vreg_28_2), .down(vreg_28_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_1), .sw(sw));
	wire signed[17:0] vwire_28_2;
	reg signed[17:0] vreg_28_2;
	node n28_2(.left(vreg_27_2), .right(vreg_29_2), .up(vreg_28_3), .down(vreg_28_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_2), .sw(sw));
	wire signed[17:0] vwire_28_3;
	reg signed[17:0] vreg_28_3;
	node n28_3(.left(vreg_27_3), .right(vreg_29_3), .up(vreg_28_4), .down(vreg_28_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_3), .sw(sw));
	wire signed[17:0] vwire_28_4;
	reg signed[17:0] vreg_28_4;
	node n28_4(.left(vreg_27_4), .right(vreg_29_4), .up(vreg_28_5), .down(vreg_28_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_4), .sw(sw));
	wire signed[17:0] vwire_28_5;
	reg signed[17:0] vreg_28_5;
	node n28_5(.left(vreg_27_5), .right(vreg_29_5), .up(vreg_28_6), .down(vreg_28_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_5), .sw(sw));
	wire signed[17:0] vwire_28_6;
	reg signed[17:0] vreg_28_6;
	node n28_6(.left(vreg_27_6), .right(vreg_29_6), .up(vreg_28_7), .down(vreg_28_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_6), .sw(sw));
	wire signed[17:0] vwire_28_7;
	reg signed[17:0] vreg_28_7;
	node n28_7(.left(vreg_27_7), .right(vreg_29_7), .up(vreg_28_8), .down(vreg_28_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_7), .sw(sw));
	wire signed[17:0] vwire_28_8;
	reg signed[17:0] vreg_28_8;
	node n28_8(.left(vreg_27_8), .right(vreg_29_8), .up(vreg_28_9), .down(vreg_28_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_8), .sw(sw));
	wire signed[17:0] vwire_28_9;
	reg signed[17:0] vreg_28_9;
	node n28_9(.left(vreg_27_9), .right(vreg_29_9), .up(vreg_28_10), .down(vreg_28_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_9), .sw(sw));
	wire signed[17:0] vwire_28_10;
	reg signed[17:0] vreg_28_10;
	node n28_10(.left(vreg_27_10), .right(vreg_29_10), .up(vreg_28_11), .down(vreg_28_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_10), .sw(sw));
	wire signed[17:0] vwire_28_11;
	reg signed[17:0] vreg_28_11;
	node n28_11(.left(vreg_27_11), .right(vreg_29_11), .up(vreg_28_12), .down(vreg_28_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_11), .sw(sw));
	wire signed[17:0] vwire_28_12;
	reg signed[17:0] vreg_28_12;
	node n28_12(.left(vreg_27_12), .right(vreg_29_12), .up(vreg_28_13), .down(vreg_28_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_12), .sw(sw));
	wire signed[17:0] vwire_28_13;
	reg signed[17:0] vreg_28_13;
	node n28_13(.left(vreg_27_13), .right(vreg_29_13), .up(vreg_28_14), .down(vreg_28_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_13), .sw(sw));
	wire signed[17:0] vwire_28_14;
	reg signed[17:0] vreg_28_14;
	node n28_14(.left(vreg_27_14), .right(vreg_29_14), .up(vreg_28_15), .down(vreg_28_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_14), .sw(sw));
	wire signed[17:0] vwire_28_15;
	reg signed[17:0] vreg_28_15;
	node n28_15(.left(vreg_27_15), .right(vreg_29_15), .up(vreg_28_16), .down(vreg_28_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_15), .sw(sw));
	wire signed[17:0] vwire_28_16;
	reg signed[17:0] vreg_28_16;
	node n28_16(.left(vreg_27_16), .right(vreg_29_16), .up(vreg_28_17), .down(vreg_28_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_16), .sw(sw));
	wire signed[17:0] vwire_28_17;
	reg signed[17:0] vreg_28_17;
	node n28_17(.left(vreg_27_17), .right(vreg_29_17), .up(vreg_28_18), .down(vreg_28_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_17), .sw(sw));
	wire signed[17:0] vwire_28_18;
	reg signed[17:0] vreg_28_18;
	node n28_18(.left(vreg_27_18), .right(vreg_29_18), .up(vreg_28_19), .down(vreg_28_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_18), .sw(sw));
	wire signed[17:0] vwire_28_19;
	reg signed[17:0] vreg_28_19;
	node n28_19(.left(vreg_27_19), .right(vreg_29_19), .up(vreg_28_20), .down(vreg_28_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_19), .sw(sw));
	wire signed[17:0] vwire_28_20;
	reg signed[17:0] vreg_28_20;
	node n28_20(.left(vreg_27_20), .right(vreg_29_20), .up(vreg_28_21), .down(vreg_28_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_20), .sw(sw));
	wire signed[17:0] vwire_28_21;
	reg signed[17:0] vreg_28_21;
	node n28_21(.left(vreg_27_21), .right(vreg_29_21), .up(vreg_28_22), .down(vreg_28_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_21), .sw(sw));
	wire signed[17:0] vwire_28_22;
	reg signed[17:0] vreg_28_22;
	node n28_22(.left(vreg_27_22), .right(vreg_29_22), .up(vreg_28_23), .down(vreg_28_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_22), .sw(sw));
	wire signed[17:0] vwire_28_23;
	reg signed[17:0] vreg_28_23;
	node n28_23(.left(vreg_27_23), .right(vreg_29_23), .up(vreg_28_24), .down(vreg_28_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_23), .sw(sw));
	wire signed[17:0] vwire_28_24;
	reg signed[17:0] vreg_28_24;
	node n28_24(.left(vreg_27_24), .right(vreg_29_24), .up(vreg_28_25), .down(vreg_28_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_24), .sw(sw));
	wire signed[17:0] vwire_28_25;
	reg signed[17:0] vreg_28_25;
	node n28_25(.left(vreg_27_25), .right(vreg_29_25), .up(vreg_28_26), .down(vreg_28_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_25), .sw(sw));
	wire signed[17:0] vwire_28_26;
	reg signed[17:0] vreg_28_26;
	node n28_26(.left(vreg_27_26), .right(vreg_29_26), .up(vreg_28_27), .down(vreg_28_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_26), .sw(sw));
	wire signed[17:0] vwire_28_27;
	reg signed[17:0] vreg_28_27;
	node n28_27(.left(vreg_27_27), .right(vreg_29_27), .up(vreg_28_28), .down(vreg_28_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_27), .sw(sw));
	wire signed[17:0] vwire_28_28;
	reg signed[17:0] vreg_28_28;
	node n28_28(.left(vreg_27_28), .right(vreg_29_28), .up(vreg_28_29), .down(vreg_28_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_28), .sw(sw));
	wire signed[17:0] vwire_28_29;
	reg signed[17:0] vreg_28_29;
	node n28_29(.left(vreg_27_29), .right(vreg_29_29), .up(vreg_28_30), .down(vreg_28_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_29), .sw(sw));
	wire signed[17:0] vwire_28_30;
	reg signed[17:0] vreg_28_30;
	node n28_30(.left(vreg_27_30), .right(vreg_29_30), .up(vreg_28_31), .down(vreg_28_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_30), .sw(sw));
	wire signed[17:0] vwire_28_31;
	reg signed[17:0] vreg_28_31;
	node n28_31(.left(vreg_27_31), .right(vreg_29_31), .up(vreg_28_32), .down(vreg_28_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_31), .sw(sw));
	wire signed[17:0] vwire_28_32;
	reg signed[17:0] vreg_28_32;
	node n28_32(.left(vreg_27_32), .right(vreg_29_32), .up(vreg_28_33), .down(vreg_28_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_32), .sw(sw));
	wire signed[17:0] vwire_28_33;
	reg signed[17:0] vreg_28_33;
	node n28_33(.left(vreg_27_33), .right(vreg_29_33), .up(vreg_28_34), .down(vreg_28_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_33), .sw(sw));
	wire signed[17:0] vwire_28_34;
	reg signed[17:0] vreg_28_34;
	node n28_34(.left(vreg_27_34), .right(vreg_29_34), .up(vreg_28_35), .down(vreg_28_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_34), .sw(sw));
	wire signed[17:0] vwire_28_35;
	reg signed[17:0] vreg_28_35;
	node n28_35(.left(vreg_27_35), .right(vreg_29_35), .up(vreg_28_36), .down(vreg_28_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_35), .sw(sw));
	wire signed[17:0] vwire_28_36;
	reg signed[17:0] vreg_28_36;
	node n28_36(.left(vreg_27_36), .right(vreg_29_36), .up(vreg_28_37), .down(vreg_28_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_36), .sw(sw));
	wire signed[17:0] vwire_28_37;
	reg signed[17:0] vreg_28_37;
	node n28_37(.left(vreg_27_37), .right(vreg_29_37), .up(vreg_28_38), .down(vreg_28_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_37), .sw(sw));
	wire signed[17:0] vwire_28_38;
	reg signed[17:0] vreg_28_38;
	node n28_38(.left(vreg_27_38), .right(vreg_29_38), .up(vreg_28_39), .down(vreg_28_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_38), .sw(sw));
	wire signed[17:0] vwire_28_39;
	reg signed[17:0] vreg_28_39;
	node n28_39(.left(vreg_27_39), .right(vreg_29_39), .up(vreg_28_40), .down(vreg_28_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_39), .sw(sw));
	wire signed[17:0] vwire_28_40;
	reg signed[17:0] vreg_28_40;
	node n28_40(.left(vreg_27_40), .right(vreg_29_40), .up(vreg_28_41), .down(vreg_28_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_40), .sw(sw));
	wire signed[17:0] vwire_28_41;
	reg signed[17:0] vreg_28_41;
	node n28_41(.left(vreg_27_41), .right(vreg_29_41), .up(vreg_28_42), .down(vreg_28_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_41), .sw(sw));
	wire signed[17:0] vwire_28_42;
	reg signed[17:0] vreg_28_42;
	node n28_42(.left(vreg_27_42), .right(vreg_29_42), .up(vreg_28_43), .down(vreg_28_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_42), .sw(sw));
	wire signed[17:0] vwire_28_43;
	reg signed[17:0] vreg_28_43;
	node n28_43(.left(vreg_27_43), .right(vreg_29_43), .up(vreg_28_44), .down(vreg_28_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_43), .sw(sw));
	wire signed[17:0] vwire_28_44;
	reg signed[17:0] vreg_28_44;
	node n28_44(.left(vreg_27_44), .right(vreg_29_44), .up(vreg_28_45), .down(vreg_28_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_44), .sw(sw));
	wire signed[17:0] vwire_28_45;
	reg signed[17:0] vreg_28_45;
	node n28_45(.left(vreg_27_45), .right(vreg_29_45), .up(vreg_28_46), .down(vreg_28_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_45), .sw(sw));
	wire signed[17:0] vwire_28_46;
	reg signed[17:0] vreg_28_46;
	node n28_46(.left(vreg_27_46), .right(vreg_29_46), .up(vreg_28_47), .down(vreg_28_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_46), .sw(sw));
	wire signed[17:0] vwire_28_47;
	reg signed[17:0] vreg_28_47;
	node n28_47(.left(vreg_27_47), .right(vreg_29_47), .up(vreg_28_48), .down(vreg_28_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_47), .sw(sw));
	wire signed[17:0] vwire_28_48;
	reg signed[17:0] vreg_28_48;
	node n28_48(.left(vreg_27_48), .right(vreg_29_48), .up(vreg_28_49), .down(vreg_28_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_48), .sw(sw));
	wire signed[17:0] vwire_28_49;
	reg signed[17:0] vreg_28_49;
	node n28_49(.left(vreg_27_49), .right(vreg_29_49), .up(18'b0), .down(vreg_28_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_28_49), .sw(sw));
	wire signed[17:0] vwire_29_0;
	reg signed[17:0] vreg_29_0;
	node n29_0(.left(vreg_28_0), .right(vreg_30_0), .up(vreg_29_1), .down(vreg_29_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_0), .sw(sw));
	wire signed[17:0] vwire_29_1;
	reg signed[17:0] vreg_29_1;
	node n29_1(.left(vreg_28_1), .right(vreg_30_1), .up(vreg_29_2), .down(vreg_29_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_1), .sw(sw));
	wire signed[17:0] vwire_29_2;
	reg signed[17:0] vreg_29_2;
	node n29_2(.left(vreg_28_2), .right(vreg_30_2), .up(vreg_29_3), .down(vreg_29_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_2), .sw(sw));
	wire signed[17:0] vwire_29_3;
	reg signed[17:0] vreg_29_3;
	node n29_3(.left(vreg_28_3), .right(vreg_30_3), .up(vreg_29_4), .down(vreg_29_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_3), .sw(sw));
	wire signed[17:0] vwire_29_4;
	reg signed[17:0] vreg_29_4;
	node n29_4(.left(vreg_28_4), .right(vreg_30_4), .up(vreg_29_5), .down(vreg_29_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_4), .sw(sw));
	wire signed[17:0] vwire_29_5;
	reg signed[17:0] vreg_29_5;
	node n29_5(.left(vreg_28_5), .right(vreg_30_5), .up(vreg_29_6), .down(vreg_29_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_5), .sw(sw));
	wire signed[17:0] vwire_29_6;
	reg signed[17:0] vreg_29_6;
	node n29_6(.left(vreg_28_6), .right(vreg_30_6), .up(vreg_29_7), .down(vreg_29_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_6), .sw(sw));
	wire signed[17:0] vwire_29_7;
	reg signed[17:0] vreg_29_7;
	node n29_7(.left(vreg_28_7), .right(vreg_30_7), .up(vreg_29_8), .down(vreg_29_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_7), .sw(sw));
	wire signed[17:0] vwire_29_8;
	reg signed[17:0] vreg_29_8;
	node n29_8(.left(vreg_28_8), .right(vreg_30_8), .up(vreg_29_9), .down(vreg_29_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_8), .sw(sw));
	wire signed[17:0] vwire_29_9;
	reg signed[17:0] vreg_29_9;
	node n29_9(.left(vreg_28_9), .right(vreg_30_9), .up(vreg_29_10), .down(vreg_29_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_9), .sw(sw));
	wire signed[17:0] vwire_29_10;
	reg signed[17:0] vreg_29_10;
	node n29_10(.left(vreg_28_10), .right(vreg_30_10), .up(vreg_29_11), .down(vreg_29_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_10), .sw(sw));
	wire signed[17:0] vwire_29_11;
	reg signed[17:0] vreg_29_11;
	node n29_11(.left(vreg_28_11), .right(vreg_30_11), .up(vreg_29_12), .down(vreg_29_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_11), .sw(sw));
	wire signed[17:0] vwire_29_12;
	reg signed[17:0] vreg_29_12;
	node n29_12(.left(vreg_28_12), .right(vreg_30_12), .up(vreg_29_13), .down(vreg_29_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_12), .sw(sw));
	wire signed[17:0] vwire_29_13;
	reg signed[17:0] vreg_29_13;
	node n29_13(.left(vreg_28_13), .right(vreg_30_13), .up(vreg_29_14), .down(vreg_29_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_13), .sw(sw));
	wire signed[17:0] vwire_29_14;
	reg signed[17:0] vreg_29_14;
	node n29_14(.left(vreg_28_14), .right(vreg_30_14), .up(vreg_29_15), .down(vreg_29_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_14), .sw(sw));
	wire signed[17:0] vwire_29_15;
	reg signed[17:0] vreg_29_15;
	node n29_15(.left(vreg_28_15), .right(vreg_30_15), .up(vreg_29_16), .down(vreg_29_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_15), .sw(sw));
	wire signed[17:0] vwire_29_16;
	reg signed[17:0] vreg_29_16;
	node n29_16(.left(vreg_28_16), .right(vreg_30_16), .up(vreg_29_17), .down(vreg_29_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_16), .sw(sw));
	wire signed[17:0] vwire_29_17;
	reg signed[17:0] vreg_29_17;
	node n29_17(.left(vreg_28_17), .right(vreg_30_17), .up(vreg_29_18), .down(vreg_29_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_17), .sw(sw));
	wire signed[17:0] vwire_29_18;
	reg signed[17:0] vreg_29_18;
	node n29_18(.left(vreg_28_18), .right(vreg_30_18), .up(vreg_29_19), .down(vreg_29_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_18), .sw(sw));
	wire signed[17:0] vwire_29_19;
	reg signed[17:0] vreg_29_19;
	node n29_19(.left(vreg_28_19), .right(vreg_30_19), .up(vreg_29_20), .down(vreg_29_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_19), .sw(sw));
	wire signed[17:0] vwire_29_20;
	reg signed[17:0] vreg_29_20;
	node n29_20(.left(vreg_28_20), .right(vreg_30_20), .up(vreg_29_21), .down(vreg_29_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_20), .sw(sw));
	wire signed[17:0] vwire_29_21;
	reg signed[17:0] vreg_29_21;
	node n29_21(.left(vreg_28_21), .right(vreg_30_21), .up(vreg_29_22), .down(vreg_29_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_21), .sw(sw));
	wire signed[17:0] vwire_29_22;
	reg signed[17:0] vreg_29_22;
	node n29_22(.left(vreg_28_22), .right(vreg_30_22), .up(vreg_29_23), .down(vreg_29_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_22), .sw(sw));
	wire signed[17:0] vwire_29_23;
	reg signed[17:0] vreg_29_23;
	node n29_23(.left(vreg_28_23), .right(vreg_30_23), .up(vreg_29_24), .down(vreg_29_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_23), .sw(sw));
	wire signed[17:0] vwire_29_24;
	reg signed[17:0] vreg_29_24;
	node n29_24(.left(vreg_28_24), .right(vreg_30_24), .up(vreg_29_25), .down(vreg_29_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_24), .sw(sw));
	wire signed[17:0] vwire_29_25;
	reg signed[17:0] vreg_29_25;
	node n29_25(.left(vreg_28_25), .right(vreg_30_25), .up(vreg_29_26), .down(vreg_29_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_25), .sw(sw));
	wire signed[17:0] vwire_29_26;
	reg signed[17:0] vreg_29_26;
	node n29_26(.left(vreg_28_26), .right(vreg_30_26), .up(vreg_29_27), .down(vreg_29_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_26), .sw(sw));
	wire signed[17:0] vwire_29_27;
	reg signed[17:0] vreg_29_27;
	node n29_27(.left(vreg_28_27), .right(vreg_30_27), .up(vreg_29_28), .down(vreg_29_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_27), .sw(sw));
	wire signed[17:0] vwire_29_28;
	reg signed[17:0] vreg_29_28;
	node n29_28(.left(vreg_28_28), .right(vreg_30_28), .up(vreg_29_29), .down(vreg_29_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_28), .sw(sw));
	wire signed[17:0] vwire_29_29;
	reg signed[17:0] vreg_29_29;
	node n29_29(.left(vreg_28_29), .right(vreg_30_29), .up(vreg_29_30), .down(vreg_29_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_29), .sw(sw));
	wire signed[17:0] vwire_29_30;
	reg signed[17:0] vreg_29_30;
	node n29_30(.left(vreg_28_30), .right(vreg_30_30), .up(vreg_29_31), .down(vreg_29_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_30), .sw(sw));
	wire signed[17:0] vwire_29_31;
	reg signed[17:0] vreg_29_31;
	node n29_31(.left(vreg_28_31), .right(vreg_30_31), .up(vreg_29_32), .down(vreg_29_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_31), .sw(sw));
	wire signed[17:0] vwire_29_32;
	reg signed[17:0] vreg_29_32;
	node n29_32(.left(vreg_28_32), .right(vreg_30_32), .up(vreg_29_33), .down(vreg_29_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_32), .sw(sw));
	wire signed[17:0] vwire_29_33;
	reg signed[17:0] vreg_29_33;
	node n29_33(.left(vreg_28_33), .right(vreg_30_33), .up(vreg_29_34), .down(vreg_29_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_33), .sw(sw));
	wire signed[17:0] vwire_29_34;
	reg signed[17:0] vreg_29_34;
	node n29_34(.left(vreg_28_34), .right(vreg_30_34), .up(vreg_29_35), .down(vreg_29_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_34), .sw(sw));
	wire signed[17:0] vwire_29_35;
	reg signed[17:0] vreg_29_35;
	node n29_35(.left(vreg_28_35), .right(vreg_30_35), .up(vreg_29_36), .down(vreg_29_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_35), .sw(sw));
	wire signed[17:0] vwire_29_36;
	reg signed[17:0] vreg_29_36;
	node n29_36(.left(vreg_28_36), .right(vreg_30_36), .up(vreg_29_37), .down(vreg_29_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_36), .sw(sw));
	wire signed[17:0] vwire_29_37;
	reg signed[17:0] vreg_29_37;
	node n29_37(.left(vreg_28_37), .right(vreg_30_37), .up(vreg_29_38), .down(vreg_29_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_37), .sw(sw));
	wire signed[17:0] vwire_29_38;
	reg signed[17:0] vreg_29_38;
	node n29_38(.left(vreg_28_38), .right(vreg_30_38), .up(vreg_29_39), .down(vreg_29_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_38), .sw(sw));
	wire signed[17:0] vwire_29_39;
	reg signed[17:0] vreg_29_39;
	node n29_39(.left(vreg_28_39), .right(vreg_30_39), .up(vreg_29_40), .down(vreg_29_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_39), .sw(sw));
	wire signed[17:0] vwire_29_40;
	reg signed[17:0] vreg_29_40;
	node n29_40(.left(vreg_28_40), .right(vreg_30_40), .up(vreg_29_41), .down(vreg_29_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_40), .sw(sw));
	wire signed[17:0] vwire_29_41;
	reg signed[17:0] vreg_29_41;
	node n29_41(.left(vreg_28_41), .right(vreg_30_41), .up(vreg_29_42), .down(vreg_29_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_41), .sw(sw));
	wire signed[17:0] vwire_29_42;
	reg signed[17:0] vreg_29_42;
	node n29_42(.left(vreg_28_42), .right(vreg_30_42), .up(vreg_29_43), .down(vreg_29_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_42), .sw(sw));
	wire signed[17:0] vwire_29_43;
	reg signed[17:0] vreg_29_43;
	node n29_43(.left(vreg_28_43), .right(vreg_30_43), .up(vreg_29_44), .down(vreg_29_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_43), .sw(sw));
	wire signed[17:0] vwire_29_44;
	reg signed[17:0] vreg_29_44;
	node n29_44(.left(vreg_28_44), .right(vreg_30_44), .up(vreg_29_45), .down(vreg_29_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_44), .sw(sw));
	wire signed[17:0] vwire_29_45;
	reg signed[17:0] vreg_29_45;
	node n29_45(.left(vreg_28_45), .right(vreg_30_45), .up(vreg_29_46), .down(vreg_29_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_45), .sw(sw));
	wire signed[17:0] vwire_29_46;
	reg signed[17:0] vreg_29_46;
	node n29_46(.left(vreg_28_46), .right(vreg_30_46), .up(vreg_29_47), .down(vreg_29_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_46), .sw(sw));
	wire signed[17:0] vwire_29_47;
	reg signed[17:0] vreg_29_47;
	node n29_47(.left(vreg_28_47), .right(vreg_30_47), .up(vreg_29_48), .down(vreg_29_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_47), .sw(sw));
	wire signed[17:0] vwire_29_48;
	reg signed[17:0] vreg_29_48;
	node n29_48(.left(vreg_28_48), .right(vreg_30_48), .up(vreg_29_49), .down(vreg_29_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_48), .sw(sw));
	wire signed[17:0] vwire_29_49;
	reg signed[17:0] vreg_29_49;
	node n29_49(.left(vreg_28_49), .right(vreg_30_49), .up(18'b0), .down(vreg_29_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_29_49), .sw(sw));
	wire signed[17:0] vwire_30_0;
	reg signed[17:0] vreg_30_0;
	node n30_0(.left(vreg_29_0), .right(vreg_31_0), .up(vreg_30_1), .down(vreg_30_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_0), .sw(sw));
	wire signed[17:0] vwire_30_1;
	reg signed[17:0] vreg_30_1;
	node n30_1(.left(vreg_29_1), .right(vreg_31_1), .up(vreg_30_2), .down(vreg_30_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_1), .sw(sw));
	wire signed[17:0] vwire_30_2;
	reg signed[17:0] vreg_30_2;
	node n30_2(.left(vreg_29_2), .right(vreg_31_2), .up(vreg_30_3), .down(vreg_30_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_2), .sw(sw));
	wire signed[17:0] vwire_30_3;
	reg signed[17:0] vreg_30_3;
	node n30_3(.left(vreg_29_3), .right(vreg_31_3), .up(vreg_30_4), .down(vreg_30_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_3), .sw(sw));
	wire signed[17:0] vwire_30_4;
	reg signed[17:0] vreg_30_4;
	node n30_4(.left(vreg_29_4), .right(vreg_31_4), .up(vreg_30_5), .down(vreg_30_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_4), .sw(sw));
	wire signed[17:0] vwire_30_5;
	reg signed[17:0] vreg_30_5;
	node n30_5(.left(vreg_29_5), .right(vreg_31_5), .up(vreg_30_6), .down(vreg_30_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_5), .sw(sw));
	wire signed[17:0] vwire_30_6;
	reg signed[17:0] vreg_30_6;
	node n30_6(.left(vreg_29_6), .right(vreg_31_6), .up(vreg_30_7), .down(vreg_30_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_6), .sw(sw));
	wire signed[17:0] vwire_30_7;
	reg signed[17:0] vreg_30_7;
	node n30_7(.left(vreg_29_7), .right(vreg_31_7), .up(vreg_30_8), .down(vreg_30_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_7), .sw(sw));
	wire signed[17:0] vwire_30_8;
	reg signed[17:0] vreg_30_8;
	node n30_8(.left(vreg_29_8), .right(vreg_31_8), .up(vreg_30_9), .down(vreg_30_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_8), .sw(sw));
	wire signed[17:0] vwire_30_9;
	reg signed[17:0] vreg_30_9;
	node n30_9(.left(vreg_29_9), .right(vreg_31_9), .up(vreg_30_10), .down(vreg_30_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_9), .sw(sw));
	wire signed[17:0] vwire_30_10;
	reg signed[17:0] vreg_30_10;
	node n30_10(.left(vreg_29_10), .right(vreg_31_10), .up(vreg_30_11), .down(vreg_30_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_10), .sw(sw));
	wire signed[17:0] vwire_30_11;
	reg signed[17:0] vreg_30_11;
	node n30_11(.left(vreg_29_11), .right(vreg_31_11), .up(vreg_30_12), .down(vreg_30_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_11), .sw(sw));
	wire signed[17:0] vwire_30_12;
	reg signed[17:0] vreg_30_12;
	node n30_12(.left(vreg_29_12), .right(vreg_31_12), .up(vreg_30_13), .down(vreg_30_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_12), .sw(sw));
	wire signed[17:0] vwire_30_13;
	reg signed[17:0] vreg_30_13;
	node n30_13(.left(vreg_29_13), .right(vreg_31_13), .up(vreg_30_14), .down(vreg_30_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_13), .sw(sw));
	wire signed[17:0] vwire_30_14;
	reg signed[17:0] vreg_30_14;
	node n30_14(.left(vreg_29_14), .right(vreg_31_14), .up(vreg_30_15), .down(vreg_30_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_14), .sw(sw));
	wire signed[17:0] vwire_30_15;
	reg signed[17:0] vreg_30_15;
	node n30_15(.left(vreg_29_15), .right(vreg_31_15), .up(vreg_30_16), .down(vreg_30_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_15), .sw(sw));
	wire signed[17:0] vwire_30_16;
	reg signed[17:0] vreg_30_16;
	node n30_16(.left(vreg_29_16), .right(vreg_31_16), .up(vreg_30_17), .down(vreg_30_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_16), .sw(sw));
	wire signed[17:0] vwire_30_17;
	reg signed[17:0] vreg_30_17;
	node n30_17(.left(vreg_29_17), .right(vreg_31_17), .up(vreg_30_18), .down(vreg_30_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_17), .sw(sw));
	wire signed[17:0] vwire_30_18;
	reg signed[17:0] vreg_30_18;
	node n30_18(.left(vreg_29_18), .right(vreg_31_18), .up(vreg_30_19), .down(vreg_30_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_18), .sw(sw));
	wire signed[17:0] vwire_30_19;
	reg signed[17:0] vreg_30_19;
	node n30_19(.left(vreg_29_19), .right(vreg_31_19), .up(vreg_30_20), .down(vreg_30_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_19), .sw(sw));
	wire signed[17:0] vwire_30_20;
	reg signed[17:0] vreg_30_20;
	node n30_20(.left(vreg_29_20), .right(vreg_31_20), .up(vreg_30_21), .down(vreg_30_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_20), .sw(sw));
	wire signed[17:0] vwire_30_21;
	reg signed[17:0] vreg_30_21;
	node n30_21(.left(vreg_29_21), .right(vreg_31_21), .up(vreg_30_22), .down(vreg_30_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_21), .sw(sw));
	wire signed[17:0] vwire_30_22;
	reg signed[17:0] vreg_30_22;
	node n30_22(.left(vreg_29_22), .right(vreg_31_22), .up(vreg_30_23), .down(vreg_30_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_22), .sw(sw));
	wire signed[17:0] vwire_30_23;
	reg signed[17:0] vreg_30_23;
	node n30_23(.left(vreg_29_23), .right(vreg_31_23), .up(vreg_30_24), .down(vreg_30_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_23), .sw(sw));
	wire signed[17:0] vwire_30_24;
	reg signed[17:0] vreg_30_24;
	node n30_24(.left(vreg_29_24), .right(vreg_31_24), .up(vreg_30_25), .down(vreg_30_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_24), .sw(sw));
	wire signed[17:0] vwire_30_25;
	reg signed[17:0] vreg_30_25;
	node n30_25(.left(vreg_29_25), .right(vreg_31_25), .up(vreg_30_26), .down(vreg_30_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_25), .sw(sw));
	wire signed[17:0] vwire_30_26;
	reg signed[17:0] vreg_30_26;
	node n30_26(.left(vreg_29_26), .right(vreg_31_26), .up(vreg_30_27), .down(vreg_30_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_26), .sw(sw));
	wire signed[17:0] vwire_30_27;
	reg signed[17:0] vreg_30_27;
	node n30_27(.left(vreg_29_27), .right(vreg_31_27), .up(vreg_30_28), .down(vreg_30_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_27), .sw(sw));
	wire signed[17:0] vwire_30_28;
	reg signed[17:0] vreg_30_28;
	node n30_28(.left(vreg_29_28), .right(vreg_31_28), .up(vreg_30_29), .down(vreg_30_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_28), .sw(sw));
	wire signed[17:0] vwire_30_29;
	reg signed[17:0] vreg_30_29;
	node n30_29(.left(vreg_29_29), .right(vreg_31_29), .up(vreg_30_30), .down(vreg_30_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_29), .sw(sw));
	wire signed[17:0] vwire_30_30;
	reg signed[17:0] vreg_30_30;
	node n30_30(.left(vreg_29_30), .right(vreg_31_30), .up(vreg_30_31), .down(vreg_30_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_30), .sw(sw));
	wire signed[17:0] vwire_30_31;
	reg signed[17:0] vreg_30_31;
	node n30_31(.left(vreg_29_31), .right(vreg_31_31), .up(vreg_30_32), .down(vreg_30_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_31), .sw(sw));
	wire signed[17:0] vwire_30_32;
	reg signed[17:0] vreg_30_32;
	node n30_32(.left(vreg_29_32), .right(vreg_31_32), .up(vreg_30_33), .down(vreg_30_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_32), .sw(sw));
	wire signed[17:0] vwire_30_33;
	reg signed[17:0] vreg_30_33;
	node n30_33(.left(vreg_29_33), .right(vreg_31_33), .up(vreg_30_34), .down(vreg_30_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_33), .sw(sw));
	wire signed[17:0] vwire_30_34;
	reg signed[17:0] vreg_30_34;
	node n30_34(.left(vreg_29_34), .right(vreg_31_34), .up(vreg_30_35), .down(vreg_30_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_34), .sw(sw));
	wire signed[17:0] vwire_30_35;
	reg signed[17:0] vreg_30_35;
	node n30_35(.left(vreg_29_35), .right(vreg_31_35), .up(vreg_30_36), .down(vreg_30_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_35), .sw(sw));
	wire signed[17:0] vwire_30_36;
	reg signed[17:0] vreg_30_36;
	node n30_36(.left(vreg_29_36), .right(vreg_31_36), .up(vreg_30_37), .down(vreg_30_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_36), .sw(sw));
	wire signed[17:0] vwire_30_37;
	reg signed[17:0] vreg_30_37;
	node n30_37(.left(vreg_29_37), .right(vreg_31_37), .up(vreg_30_38), .down(vreg_30_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_37), .sw(sw));
	wire signed[17:0] vwire_30_38;
	reg signed[17:0] vreg_30_38;
	node n30_38(.left(vreg_29_38), .right(vreg_31_38), .up(vreg_30_39), .down(vreg_30_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_38), .sw(sw));
	wire signed[17:0] vwire_30_39;
	reg signed[17:0] vreg_30_39;
	node n30_39(.left(vreg_29_39), .right(vreg_31_39), .up(vreg_30_40), .down(vreg_30_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_39), .sw(sw));
	wire signed[17:0] vwire_30_40;
	reg signed[17:0] vreg_30_40;
	node n30_40(.left(vreg_29_40), .right(vreg_31_40), .up(vreg_30_41), .down(vreg_30_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_40), .sw(sw));
	wire signed[17:0] vwire_30_41;
	reg signed[17:0] vreg_30_41;
	node n30_41(.left(vreg_29_41), .right(vreg_31_41), .up(vreg_30_42), .down(vreg_30_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_41), .sw(sw));
	wire signed[17:0] vwire_30_42;
	reg signed[17:0] vreg_30_42;
	node n30_42(.left(vreg_29_42), .right(vreg_31_42), .up(vreg_30_43), .down(vreg_30_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_42), .sw(sw));
	wire signed[17:0] vwire_30_43;
	reg signed[17:0] vreg_30_43;
	node n30_43(.left(vreg_29_43), .right(vreg_31_43), .up(vreg_30_44), .down(vreg_30_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_43), .sw(sw));
	wire signed[17:0] vwire_30_44;
	reg signed[17:0] vreg_30_44;
	node n30_44(.left(vreg_29_44), .right(vreg_31_44), .up(vreg_30_45), .down(vreg_30_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_44), .sw(sw));
	wire signed[17:0] vwire_30_45;
	reg signed[17:0] vreg_30_45;
	node n30_45(.left(vreg_29_45), .right(vreg_31_45), .up(vreg_30_46), .down(vreg_30_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_45), .sw(sw));
	wire signed[17:0] vwire_30_46;
	reg signed[17:0] vreg_30_46;
	node n30_46(.left(vreg_29_46), .right(vreg_31_46), .up(vreg_30_47), .down(vreg_30_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_46), .sw(sw));
	wire signed[17:0] vwire_30_47;
	reg signed[17:0] vreg_30_47;
	node n30_47(.left(vreg_29_47), .right(vreg_31_47), .up(vreg_30_48), .down(vreg_30_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_47), .sw(sw));
	wire signed[17:0] vwire_30_48;
	reg signed[17:0] vreg_30_48;
	node n30_48(.left(vreg_29_48), .right(vreg_31_48), .up(vreg_30_49), .down(vreg_30_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_48), .sw(sw));
	wire signed[17:0] vwire_30_49;
	reg signed[17:0] vreg_30_49;
	node n30_49(.left(vreg_29_49), .right(vreg_31_49), .up(18'b0), .down(vreg_30_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_30_49), .sw(sw));
	wire signed[17:0] vwire_31_0;
	reg signed[17:0] vreg_31_0;
	node n31_0(.left(vreg_30_0), .right(vreg_32_0), .up(vreg_31_1), .down(vreg_31_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_0), .sw(sw));
	wire signed[17:0] vwire_31_1;
	reg signed[17:0] vreg_31_1;
	node n31_1(.left(vreg_30_1), .right(vreg_32_1), .up(vreg_31_2), .down(vreg_31_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_1), .sw(sw));
	wire signed[17:0] vwire_31_2;
	reg signed[17:0] vreg_31_2;
	node n31_2(.left(vreg_30_2), .right(vreg_32_2), .up(vreg_31_3), .down(vreg_31_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_2), .sw(sw));
	wire signed[17:0] vwire_31_3;
	reg signed[17:0] vreg_31_3;
	node n31_3(.left(vreg_30_3), .right(vreg_32_3), .up(vreg_31_4), .down(vreg_31_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_3), .sw(sw));
	wire signed[17:0] vwire_31_4;
	reg signed[17:0] vreg_31_4;
	node n31_4(.left(vreg_30_4), .right(vreg_32_4), .up(vreg_31_5), .down(vreg_31_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_4), .sw(sw));
	wire signed[17:0] vwire_31_5;
	reg signed[17:0] vreg_31_5;
	node n31_5(.left(vreg_30_5), .right(vreg_32_5), .up(vreg_31_6), .down(vreg_31_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_5), .sw(sw));
	wire signed[17:0] vwire_31_6;
	reg signed[17:0] vreg_31_6;
	node n31_6(.left(vreg_30_6), .right(vreg_32_6), .up(vreg_31_7), .down(vreg_31_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_6), .sw(sw));
	wire signed[17:0] vwire_31_7;
	reg signed[17:0] vreg_31_7;
	node n31_7(.left(vreg_30_7), .right(vreg_32_7), .up(vreg_31_8), .down(vreg_31_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_7), .sw(sw));
	wire signed[17:0] vwire_31_8;
	reg signed[17:0] vreg_31_8;
	node n31_8(.left(vreg_30_8), .right(vreg_32_8), .up(vreg_31_9), .down(vreg_31_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_8), .sw(sw));
	wire signed[17:0] vwire_31_9;
	reg signed[17:0] vreg_31_9;
	node n31_9(.left(vreg_30_9), .right(vreg_32_9), .up(vreg_31_10), .down(vreg_31_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_9), .sw(sw));
	wire signed[17:0] vwire_31_10;
	reg signed[17:0] vreg_31_10;
	node n31_10(.left(vreg_30_10), .right(vreg_32_10), .up(vreg_31_11), .down(vreg_31_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_10), .sw(sw));
	wire signed[17:0] vwire_31_11;
	reg signed[17:0] vreg_31_11;
	node n31_11(.left(vreg_30_11), .right(vreg_32_11), .up(vreg_31_12), .down(vreg_31_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_11), .sw(sw));
	wire signed[17:0] vwire_31_12;
	reg signed[17:0] vreg_31_12;
	node n31_12(.left(vreg_30_12), .right(vreg_32_12), .up(vreg_31_13), .down(vreg_31_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_12), .sw(sw));
	wire signed[17:0] vwire_31_13;
	reg signed[17:0] vreg_31_13;
	node n31_13(.left(vreg_30_13), .right(vreg_32_13), .up(vreg_31_14), .down(vreg_31_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_13), .sw(sw));
	wire signed[17:0] vwire_31_14;
	reg signed[17:0] vreg_31_14;
	node n31_14(.left(vreg_30_14), .right(vreg_32_14), .up(vreg_31_15), .down(vreg_31_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_14), .sw(sw));
	wire signed[17:0] vwire_31_15;
	reg signed[17:0] vreg_31_15;
	node n31_15(.left(vreg_30_15), .right(vreg_32_15), .up(vreg_31_16), .down(vreg_31_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_15), .sw(sw));
	wire signed[17:0] vwire_31_16;
	reg signed[17:0] vreg_31_16;
	node n31_16(.left(vreg_30_16), .right(vreg_32_16), .up(vreg_31_17), .down(vreg_31_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_16), .sw(sw));
	wire signed[17:0] vwire_31_17;
	reg signed[17:0] vreg_31_17;
	node n31_17(.left(vreg_30_17), .right(vreg_32_17), .up(vreg_31_18), .down(vreg_31_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_17), .sw(sw));
	wire signed[17:0] vwire_31_18;
	reg signed[17:0] vreg_31_18;
	node n31_18(.left(vreg_30_18), .right(vreg_32_18), .up(vreg_31_19), .down(vreg_31_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_18), .sw(sw));
	wire signed[17:0] vwire_31_19;
	reg signed[17:0] vreg_31_19;
	node n31_19(.left(vreg_30_19), .right(vreg_32_19), .up(vreg_31_20), .down(vreg_31_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_19), .sw(sw));
	wire signed[17:0] vwire_31_20;
	reg signed[17:0] vreg_31_20;
	node n31_20(.left(vreg_30_20), .right(vreg_32_20), .up(vreg_31_21), .down(vreg_31_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_20), .sw(sw));
	wire signed[17:0] vwire_31_21;
	reg signed[17:0] vreg_31_21;
	node n31_21(.left(vreg_30_21), .right(vreg_32_21), .up(vreg_31_22), .down(vreg_31_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_21), .sw(sw));
	wire signed[17:0] vwire_31_22;
	reg signed[17:0] vreg_31_22;
	node n31_22(.left(vreg_30_22), .right(vreg_32_22), .up(vreg_31_23), .down(vreg_31_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_22), .sw(sw));
	wire signed[17:0] vwire_31_23;
	reg signed[17:0] vreg_31_23;
	node n31_23(.left(vreg_30_23), .right(vreg_32_23), .up(vreg_31_24), .down(vreg_31_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_23), .sw(sw));
	wire signed[17:0] vwire_31_24;
	reg signed[17:0] vreg_31_24;
	node n31_24(.left(vreg_30_24), .right(vreg_32_24), .up(vreg_31_25), .down(vreg_31_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_24), .sw(sw));
	wire signed[17:0] vwire_31_25;
	reg signed[17:0] vreg_31_25;
	node n31_25(.left(vreg_30_25), .right(vreg_32_25), .up(vreg_31_26), .down(vreg_31_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_25), .sw(sw));
	wire signed[17:0] vwire_31_26;
	reg signed[17:0] vreg_31_26;
	node n31_26(.left(vreg_30_26), .right(vreg_32_26), .up(vreg_31_27), .down(vreg_31_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_26), .sw(sw));
	wire signed[17:0] vwire_31_27;
	reg signed[17:0] vreg_31_27;
	node n31_27(.left(vreg_30_27), .right(vreg_32_27), .up(vreg_31_28), .down(vreg_31_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_27), .sw(sw));
	wire signed[17:0] vwire_31_28;
	reg signed[17:0] vreg_31_28;
	node n31_28(.left(vreg_30_28), .right(vreg_32_28), .up(vreg_31_29), .down(vreg_31_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_28), .sw(sw));
	wire signed[17:0] vwire_31_29;
	reg signed[17:0] vreg_31_29;
	node n31_29(.left(vreg_30_29), .right(vreg_32_29), .up(vreg_31_30), .down(vreg_31_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_29), .sw(sw));
	wire signed[17:0] vwire_31_30;
	reg signed[17:0] vreg_31_30;
	node n31_30(.left(vreg_30_30), .right(vreg_32_30), .up(vreg_31_31), .down(vreg_31_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_30), .sw(sw));
	wire signed[17:0] vwire_31_31;
	reg signed[17:0] vreg_31_31;
	node n31_31(.left(vreg_30_31), .right(vreg_32_31), .up(vreg_31_32), .down(vreg_31_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_31), .sw(sw));
	wire signed[17:0] vwire_31_32;
	reg signed[17:0] vreg_31_32;
	node n31_32(.left(vreg_30_32), .right(vreg_32_32), .up(vreg_31_33), .down(vreg_31_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_32), .sw(sw));
	wire signed[17:0] vwire_31_33;
	reg signed[17:0] vreg_31_33;
	node n31_33(.left(vreg_30_33), .right(vreg_32_33), .up(vreg_31_34), .down(vreg_31_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_33), .sw(sw));
	wire signed[17:0] vwire_31_34;
	reg signed[17:0] vreg_31_34;
	node n31_34(.left(vreg_30_34), .right(vreg_32_34), .up(vreg_31_35), .down(vreg_31_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_34), .sw(sw));
	wire signed[17:0] vwire_31_35;
	reg signed[17:0] vreg_31_35;
	node n31_35(.left(vreg_30_35), .right(vreg_32_35), .up(vreg_31_36), .down(vreg_31_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_35), .sw(sw));
	wire signed[17:0] vwire_31_36;
	reg signed[17:0] vreg_31_36;
	node n31_36(.left(vreg_30_36), .right(vreg_32_36), .up(vreg_31_37), .down(vreg_31_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_36), .sw(sw));
	wire signed[17:0] vwire_31_37;
	reg signed[17:0] vreg_31_37;
	node n31_37(.left(vreg_30_37), .right(vreg_32_37), .up(vreg_31_38), .down(vreg_31_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_37), .sw(sw));
	wire signed[17:0] vwire_31_38;
	reg signed[17:0] vreg_31_38;
	node n31_38(.left(vreg_30_38), .right(vreg_32_38), .up(vreg_31_39), .down(vreg_31_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_38), .sw(sw));
	wire signed[17:0] vwire_31_39;
	reg signed[17:0] vreg_31_39;
	node n31_39(.left(vreg_30_39), .right(vreg_32_39), .up(vreg_31_40), .down(vreg_31_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_39), .sw(sw));
	wire signed[17:0] vwire_31_40;
	reg signed[17:0] vreg_31_40;
	node n31_40(.left(vreg_30_40), .right(vreg_32_40), .up(vreg_31_41), .down(vreg_31_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_40), .sw(sw));
	wire signed[17:0] vwire_31_41;
	reg signed[17:0] vreg_31_41;
	node n31_41(.left(vreg_30_41), .right(vreg_32_41), .up(vreg_31_42), .down(vreg_31_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_41), .sw(sw));
	wire signed[17:0] vwire_31_42;
	reg signed[17:0] vreg_31_42;
	node n31_42(.left(vreg_30_42), .right(vreg_32_42), .up(vreg_31_43), .down(vreg_31_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_42), .sw(sw));
	wire signed[17:0] vwire_31_43;
	reg signed[17:0] vreg_31_43;
	node n31_43(.left(vreg_30_43), .right(vreg_32_43), .up(vreg_31_44), .down(vreg_31_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_43), .sw(sw));
	wire signed[17:0] vwire_31_44;
	reg signed[17:0] vreg_31_44;
	node n31_44(.left(vreg_30_44), .right(vreg_32_44), .up(vreg_31_45), .down(vreg_31_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_44), .sw(sw));
	wire signed[17:0] vwire_31_45;
	reg signed[17:0] vreg_31_45;
	node n31_45(.left(vreg_30_45), .right(vreg_32_45), .up(vreg_31_46), .down(vreg_31_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_45), .sw(sw));
	wire signed[17:0] vwire_31_46;
	reg signed[17:0] vreg_31_46;
	node n31_46(.left(vreg_30_46), .right(vreg_32_46), .up(vreg_31_47), .down(vreg_31_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_46), .sw(sw));
	wire signed[17:0] vwire_31_47;
	reg signed[17:0] vreg_31_47;
	node n31_47(.left(vreg_30_47), .right(vreg_32_47), .up(vreg_31_48), .down(vreg_31_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_47), .sw(sw));
	wire signed[17:0] vwire_31_48;
	reg signed[17:0] vreg_31_48;
	node n31_48(.left(vreg_30_48), .right(vreg_32_48), .up(vreg_31_49), .down(vreg_31_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_48), .sw(sw));
	wire signed[17:0] vwire_31_49;
	reg signed[17:0] vreg_31_49;
	node n31_49(.left(vreg_30_49), .right(vreg_32_49), .up(18'b0), .down(vreg_31_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_31_49), .sw(sw));
	wire signed[17:0] vwire_32_0;
	reg signed[17:0] vreg_32_0;
	node n32_0(.left(vreg_31_0), .right(vreg_33_0), .up(vreg_32_1), .down(vreg_32_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_0), .sw(sw));
	wire signed[17:0] vwire_32_1;
	reg signed[17:0] vreg_32_1;
	node n32_1(.left(vreg_31_1), .right(vreg_33_1), .up(vreg_32_2), .down(vreg_32_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_1), .sw(sw));
	wire signed[17:0] vwire_32_2;
	reg signed[17:0] vreg_32_2;
	node n32_2(.left(vreg_31_2), .right(vreg_33_2), .up(vreg_32_3), .down(vreg_32_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_2), .sw(sw));
	wire signed[17:0] vwire_32_3;
	reg signed[17:0] vreg_32_3;
	node n32_3(.left(vreg_31_3), .right(vreg_33_3), .up(vreg_32_4), .down(vreg_32_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_3), .sw(sw));
	wire signed[17:0] vwire_32_4;
	reg signed[17:0] vreg_32_4;
	node n32_4(.left(vreg_31_4), .right(vreg_33_4), .up(vreg_32_5), .down(vreg_32_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_4), .sw(sw));
	wire signed[17:0] vwire_32_5;
	reg signed[17:0] vreg_32_5;
	node n32_5(.left(vreg_31_5), .right(vreg_33_5), .up(vreg_32_6), .down(vreg_32_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_5), .sw(sw));
	wire signed[17:0] vwire_32_6;
	reg signed[17:0] vreg_32_6;
	node n32_6(.left(vreg_31_6), .right(vreg_33_6), .up(vreg_32_7), .down(vreg_32_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_6), .sw(sw));
	wire signed[17:0] vwire_32_7;
	reg signed[17:0] vreg_32_7;
	node n32_7(.left(vreg_31_7), .right(vreg_33_7), .up(vreg_32_8), .down(vreg_32_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_7), .sw(sw));
	wire signed[17:0] vwire_32_8;
	reg signed[17:0] vreg_32_8;
	node n32_8(.left(vreg_31_8), .right(vreg_33_8), .up(vreg_32_9), .down(vreg_32_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_8), .sw(sw));
	wire signed[17:0] vwire_32_9;
	reg signed[17:0] vreg_32_9;
	node n32_9(.left(vreg_31_9), .right(vreg_33_9), .up(vreg_32_10), .down(vreg_32_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_9), .sw(sw));
	wire signed[17:0] vwire_32_10;
	reg signed[17:0] vreg_32_10;
	node n32_10(.left(vreg_31_10), .right(vreg_33_10), .up(vreg_32_11), .down(vreg_32_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_10), .sw(sw));
	wire signed[17:0] vwire_32_11;
	reg signed[17:0] vreg_32_11;
	node n32_11(.left(vreg_31_11), .right(vreg_33_11), .up(vreg_32_12), .down(vreg_32_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_11), .sw(sw));
	wire signed[17:0] vwire_32_12;
	reg signed[17:0] vreg_32_12;
	node n32_12(.left(vreg_31_12), .right(vreg_33_12), .up(vreg_32_13), .down(vreg_32_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_12), .sw(sw));
	wire signed[17:0] vwire_32_13;
	reg signed[17:0] vreg_32_13;
	node n32_13(.left(vreg_31_13), .right(vreg_33_13), .up(vreg_32_14), .down(vreg_32_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_13), .sw(sw));
	wire signed[17:0] vwire_32_14;
	reg signed[17:0] vreg_32_14;
	node n32_14(.left(vreg_31_14), .right(vreg_33_14), .up(vreg_32_15), .down(vreg_32_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_14), .sw(sw));
	wire signed[17:0] vwire_32_15;
	reg signed[17:0] vreg_32_15;
	node n32_15(.left(vreg_31_15), .right(vreg_33_15), .up(vreg_32_16), .down(vreg_32_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_15), .sw(sw));
	wire signed[17:0] vwire_32_16;
	reg signed[17:0] vreg_32_16;
	node n32_16(.left(vreg_31_16), .right(vreg_33_16), .up(vreg_32_17), .down(vreg_32_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_16), .sw(sw));
	wire signed[17:0] vwire_32_17;
	reg signed[17:0] vreg_32_17;
	node n32_17(.left(vreg_31_17), .right(vreg_33_17), .up(vreg_32_18), .down(vreg_32_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_17), .sw(sw));
	wire signed[17:0] vwire_32_18;
	reg signed[17:0] vreg_32_18;
	node n32_18(.left(vreg_31_18), .right(vreg_33_18), .up(vreg_32_19), .down(vreg_32_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_18), .sw(sw));
	wire signed[17:0] vwire_32_19;
	reg signed[17:0] vreg_32_19;
	node n32_19(.left(vreg_31_19), .right(vreg_33_19), .up(vreg_32_20), .down(vreg_32_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_19), .sw(sw));
	wire signed[17:0] vwire_32_20;
	reg signed[17:0] vreg_32_20;
	node n32_20(.left(vreg_31_20), .right(vreg_33_20), .up(vreg_32_21), .down(vreg_32_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_20), .sw(sw));
	wire signed[17:0] vwire_32_21;
	reg signed[17:0] vreg_32_21;
	node n32_21(.left(vreg_31_21), .right(vreg_33_21), .up(vreg_32_22), .down(vreg_32_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_21), .sw(sw));
	wire signed[17:0] vwire_32_22;
	reg signed[17:0] vreg_32_22;
	node n32_22(.left(vreg_31_22), .right(vreg_33_22), .up(vreg_32_23), .down(vreg_32_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_22), .sw(sw));
	wire signed[17:0] vwire_32_23;
	reg signed[17:0] vreg_32_23;
	node n32_23(.left(vreg_31_23), .right(vreg_33_23), .up(vreg_32_24), .down(vreg_32_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_23), .sw(sw));
	wire signed[17:0] vwire_32_24;
	reg signed[17:0] vreg_32_24;
	node n32_24(.left(vreg_31_24), .right(vreg_33_24), .up(vreg_32_25), .down(vreg_32_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_24), .sw(sw));
	wire signed[17:0] vwire_32_25;
	reg signed[17:0] vreg_32_25;
	node n32_25(.left(vreg_31_25), .right(vreg_33_25), .up(vreg_32_26), .down(vreg_32_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_25), .sw(sw));
	wire signed[17:0] vwire_32_26;
	reg signed[17:0] vreg_32_26;
	node n32_26(.left(vreg_31_26), .right(vreg_33_26), .up(vreg_32_27), .down(vreg_32_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_26), .sw(sw));
	wire signed[17:0] vwire_32_27;
	reg signed[17:0] vreg_32_27;
	node n32_27(.left(vreg_31_27), .right(vreg_33_27), .up(vreg_32_28), .down(vreg_32_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_27), .sw(sw));
	wire signed[17:0] vwire_32_28;
	reg signed[17:0] vreg_32_28;
	node n32_28(.left(vreg_31_28), .right(vreg_33_28), .up(vreg_32_29), .down(vreg_32_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_28), .sw(sw));
	wire signed[17:0] vwire_32_29;
	reg signed[17:0] vreg_32_29;
	node n32_29(.left(vreg_31_29), .right(vreg_33_29), .up(vreg_32_30), .down(vreg_32_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_29), .sw(sw));
	wire signed[17:0] vwire_32_30;
	reg signed[17:0] vreg_32_30;
	node n32_30(.left(vreg_31_30), .right(vreg_33_30), .up(vreg_32_31), .down(vreg_32_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_30), .sw(sw));
	wire signed[17:0] vwire_32_31;
	reg signed[17:0] vreg_32_31;
	node n32_31(.left(vreg_31_31), .right(vreg_33_31), .up(vreg_32_32), .down(vreg_32_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_31), .sw(sw));
	wire signed[17:0] vwire_32_32;
	reg signed[17:0] vreg_32_32;
	node n32_32(.left(vreg_31_32), .right(vreg_33_32), .up(vreg_32_33), .down(vreg_32_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_32), .sw(sw));
	wire signed[17:0] vwire_32_33;
	reg signed[17:0] vreg_32_33;
	node n32_33(.left(vreg_31_33), .right(vreg_33_33), .up(vreg_32_34), .down(vreg_32_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_33), .sw(sw));
	wire signed[17:0] vwire_32_34;
	reg signed[17:0] vreg_32_34;
	node n32_34(.left(vreg_31_34), .right(vreg_33_34), .up(vreg_32_35), .down(vreg_32_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_34), .sw(sw));
	wire signed[17:0] vwire_32_35;
	reg signed[17:0] vreg_32_35;
	node n32_35(.left(vreg_31_35), .right(vreg_33_35), .up(vreg_32_36), .down(vreg_32_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_35), .sw(sw));
	wire signed[17:0] vwire_32_36;
	reg signed[17:0] vreg_32_36;
	node n32_36(.left(vreg_31_36), .right(vreg_33_36), .up(vreg_32_37), .down(vreg_32_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_36), .sw(sw));
	wire signed[17:0] vwire_32_37;
	reg signed[17:0] vreg_32_37;
	node n32_37(.left(vreg_31_37), .right(vreg_33_37), .up(vreg_32_38), .down(vreg_32_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_37), .sw(sw));
	wire signed[17:0] vwire_32_38;
	reg signed[17:0] vreg_32_38;
	node n32_38(.left(vreg_31_38), .right(vreg_33_38), .up(vreg_32_39), .down(vreg_32_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_38), .sw(sw));
	wire signed[17:0] vwire_32_39;
	reg signed[17:0] vreg_32_39;
	node n32_39(.left(vreg_31_39), .right(vreg_33_39), .up(vreg_32_40), .down(vreg_32_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_39), .sw(sw));
	wire signed[17:0] vwire_32_40;
	reg signed[17:0] vreg_32_40;
	node n32_40(.left(vreg_31_40), .right(vreg_33_40), .up(vreg_32_41), .down(vreg_32_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_40), .sw(sw));
	wire signed[17:0] vwire_32_41;
	reg signed[17:0] vreg_32_41;
	node n32_41(.left(vreg_31_41), .right(vreg_33_41), .up(vreg_32_42), .down(vreg_32_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_41), .sw(sw));
	wire signed[17:0] vwire_32_42;
	reg signed[17:0] vreg_32_42;
	node n32_42(.left(vreg_31_42), .right(vreg_33_42), .up(vreg_32_43), .down(vreg_32_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_42), .sw(sw));
	wire signed[17:0] vwire_32_43;
	reg signed[17:0] vreg_32_43;
	node n32_43(.left(vreg_31_43), .right(vreg_33_43), .up(vreg_32_44), .down(vreg_32_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_43), .sw(sw));
	wire signed[17:0] vwire_32_44;
	reg signed[17:0] vreg_32_44;
	node n32_44(.left(vreg_31_44), .right(vreg_33_44), .up(vreg_32_45), .down(vreg_32_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_44), .sw(sw));
	wire signed[17:0] vwire_32_45;
	reg signed[17:0] vreg_32_45;
	node n32_45(.left(vreg_31_45), .right(vreg_33_45), .up(vreg_32_46), .down(vreg_32_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_45), .sw(sw));
	wire signed[17:0] vwire_32_46;
	reg signed[17:0] vreg_32_46;
	node n32_46(.left(vreg_31_46), .right(vreg_33_46), .up(vreg_32_47), .down(vreg_32_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_46), .sw(sw));
	wire signed[17:0] vwire_32_47;
	reg signed[17:0] vreg_32_47;
	node n32_47(.left(vreg_31_47), .right(vreg_33_47), .up(vreg_32_48), .down(vreg_32_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_47), .sw(sw));
	wire signed[17:0] vwire_32_48;
	reg signed[17:0] vreg_32_48;
	node n32_48(.left(vreg_31_48), .right(vreg_33_48), .up(vreg_32_49), .down(vreg_32_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_48), .sw(sw));
	wire signed[17:0] vwire_32_49;
	reg signed[17:0] vreg_32_49;
	node n32_49(.left(vreg_31_49), .right(vreg_33_49), .up(18'b0), .down(vreg_32_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_32_49), .sw(sw));
	wire signed[17:0] vwire_33_0;
	reg signed[17:0] vreg_33_0;
	node n33_0(.left(vreg_32_0), .right(vreg_34_0), .up(vreg_33_1), .down(vreg_33_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_0), .sw(sw));
	wire signed[17:0] vwire_33_1;
	reg signed[17:0] vreg_33_1;
	node n33_1(.left(vreg_32_1), .right(vreg_34_1), .up(vreg_33_2), .down(vreg_33_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_1), .sw(sw));
	wire signed[17:0] vwire_33_2;
	reg signed[17:0] vreg_33_2;
	node n33_2(.left(vreg_32_2), .right(vreg_34_2), .up(vreg_33_3), .down(vreg_33_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_2), .sw(sw));
	wire signed[17:0] vwire_33_3;
	reg signed[17:0] vreg_33_3;
	node n33_3(.left(vreg_32_3), .right(vreg_34_3), .up(vreg_33_4), .down(vreg_33_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_3), .sw(sw));
	wire signed[17:0] vwire_33_4;
	reg signed[17:0] vreg_33_4;
	node n33_4(.left(vreg_32_4), .right(vreg_34_4), .up(vreg_33_5), .down(vreg_33_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_4), .sw(sw));
	wire signed[17:0] vwire_33_5;
	reg signed[17:0] vreg_33_5;
	node n33_5(.left(vreg_32_5), .right(vreg_34_5), .up(vreg_33_6), .down(vreg_33_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_5), .sw(sw));
	wire signed[17:0] vwire_33_6;
	reg signed[17:0] vreg_33_6;
	node n33_6(.left(vreg_32_6), .right(vreg_34_6), .up(vreg_33_7), .down(vreg_33_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_6), .sw(sw));
	wire signed[17:0] vwire_33_7;
	reg signed[17:0] vreg_33_7;
	node n33_7(.left(vreg_32_7), .right(vreg_34_7), .up(vreg_33_8), .down(vreg_33_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_7), .sw(sw));
	wire signed[17:0] vwire_33_8;
	reg signed[17:0] vreg_33_8;
	node n33_8(.left(vreg_32_8), .right(vreg_34_8), .up(vreg_33_9), .down(vreg_33_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_8), .sw(sw));
	wire signed[17:0] vwire_33_9;
	reg signed[17:0] vreg_33_9;
	node n33_9(.left(vreg_32_9), .right(vreg_34_9), .up(vreg_33_10), .down(vreg_33_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_9), .sw(sw));
	wire signed[17:0] vwire_33_10;
	reg signed[17:0] vreg_33_10;
	node n33_10(.left(vreg_32_10), .right(vreg_34_10), .up(vreg_33_11), .down(vreg_33_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_10), .sw(sw));
	wire signed[17:0] vwire_33_11;
	reg signed[17:0] vreg_33_11;
	node n33_11(.left(vreg_32_11), .right(vreg_34_11), .up(vreg_33_12), .down(vreg_33_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_11), .sw(sw));
	wire signed[17:0] vwire_33_12;
	reg signed[17:0] vreg_33_12;
	node n33_12(.left(vreg_32_12), .right(vreg_34_12), .up(vreg_33_13), .down(vreg_33_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_12), .sw(sw));
	wire signed[17:0] vwire_33_13;
	reg signed[17:0] vreg_33_13;
	node n33_13(.left(vreg_32_13), .right(vreg_34_13), .up(vreg_33_14), .down(vreg_33_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_13), .sw(sw));
	wire signed[17:0] vwire_33_14;
	reg signed[17:0] vreg_33_14;
	node n33_14(.left(vreg_32_14), .right(vreg_34_14), .up(vreg_33_15), .down(vreg_33_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_14), .sw(sw));
	wire signed[17:0] vwire_33_15;
	reg signed[17:0] vreg_33_15;
	node n33_15(.left(vreg_32_15), .right(vreg_34_15), .up(vreg_33_16), .down(vreg_33_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_15), .sw(sw));
	wire signed[17:0] vwire_33_16;
	reg signed[17:0] vreg_33_16;
	node n33_16(.left(vreg_32_16), .right(vreg_34_16), .up(vreg_33_17), .down(vreg_33_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_16), .sw(sw));
	wire signed[17:0] vwire_33_17;
	reg signed[17:0] vreg_33_17;
	node n33_17(.left(vreg_32_17), .right(vreg_34_17), .up(vreg_33_18), .down(vreg_33_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_17), .sw(sw));
	wire signed[17:0] vwire_33_18;
	reg signed[17:0] vreg_33_18;
	node n33_18(.left(vreg_32_18), .right(vreg_34_18), .up(vreg_33_19), .down(vreg_33_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_18), .sw(sw));
	wire signed[17:0] vwire_33_19;
	reg signed[17:0] vreg_33_19;
	node n33_19(.left(vreg_32_19), .right(vreg_34_19), .up(vreg_33_20), .down(vreg_33_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_19), .sw(sw));
	wire signed[17:0] vwire_33_20;
	reg signed[17:0] vreg_33_20;
	node n33_20(.left(vreg_32_20), .right(vreg_34_20), .up(vreg_33_21), .down(vreg_33_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_20), .sw(sw));
	wire signed[17:0] vwire_33_21;
	reg signed[17:0] vreg_33_21;
	node n33_21(.left(vreg_32_21), .right(vreg_34_21), .up(vreg_33_22), .down(vreg_33_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_21), .sw(sw));
	wire signed[17:0] vwire_33_22;
	reg signed[17:0] vreg_33_22;
	node n33_22(.left(vreg_32_22), .right(vreg_34_22), .up(vreg_33_23), .down(vreg_33_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_22), .sw(sw));
	wire signed[17:0] vwire_33_23;
	reg signed[17:0] vreg_33_23;
	node n33_23(.left(vreg_32_23), .right(vreg_34_23), .up(vreg_33_24), .down(vreg_33_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_23), .sw(sw));
	wire signed[17:0] vwire_33_24;
	reg signed[17:0] vreg_33_24;
	node n33_24(.left(vreg_32_24), .right(vreg_34_24), .up(vreg_33_25), .down(vreg_33_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_24), .sw(sw));
	wire signed[17:0] vwire_33_25;
	reg signed[17:0] vreg_33_25;
	node n33_25(.left(vreg_32_25), .right(vreg_34_25), .up(vreg_33_26), .down(vreg_33_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_25), .sw(sw));
	wire signed[17:0] vwire_33_26;
	reg signed[17:0] vreg_33_26;
	node n33_26(.left(vreg_32_26), .right(vreg_34_26), .up(vreg_33_27), .down(vreg_33_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_26), .sw(sw));
	wire signed[17:0] vwire_33_27;
	reg signed[17:0] vreg_33_27;
	node n33_27(.left(vreg_32_27), .right(vreg_34_27), .up(vreg_33_28), .down(vreg_33_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_27), .sw(sw));
	wire signed[17:0] vwire_33_28;
	reg signed[17:0] vreg_33_28;
	node n33_28(.left(vreg_32_28), .right(vreg_34_28), .up(vreg_33_29), .down(vreg_33_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_28), .sw(sw));
	wire signed[17:0] vwire_33_29;
	reg signed[17:0] vreg_33_29;
	node n33_29(.left(vreg_32_29), .right(vreg_34_29), .up(vreg_33_30), .down(vreg_33_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_29), .sw(sw));
	wire signed[17:0] vwire_33_30;
	reg signed[17:0] vreg_33_30;
	node n33_30(.left(vreg_32_30), .right(vreg_34_30), .up(vreg_33_31), .down(vreg_33_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_30), .sw(sw));
	wire signed[17:0] vwire_33_31;
	reg signed[17:0] vreg_33_31;
	node n33_31(.left(vreg_32_31), .right(vreg_34_31), .up(vreg_33_32), .down(vreg_33_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_31), .sw(sw));
	wire signed[17:0] vwire_33_32;
	reg signed[17:0] vreg_33_32;
	node n33_32(.left(vreg_32_32), .right(vreg_34_32), .up(vreg_33_33), .down(vreg_33_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_32), .sw(sw));
	wire signed[17:0] vwire_33_33;
	reg signed[17:0] vreg_33_33;
	node n33_33(.left(vreg_32_33), .right(vreg_34_33), .up(vreg_33_34), .down(vreg_33_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_33), .sw(sw));
	wire signed[17:0] vwire_33_34;
	reg signed[17:0] vreg_33_34;
	node n33_34(.left(vreg_32_34), .right(vreg_34_34), .up(vreg_33_35), .down(vreg_33_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_34), .sw(sw));
	wire signed[17:0] vwire_33_35;
	reg signed[17:0] vreg_33_35;
	node n33_35(.left(vreg_32_35), .right(vreg_34_35), .up(vreg_33_36), .down(vreg_33_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_35), .sw(sw));
	wire signed[17:0] vwire_33_36;
	reg signed[17:0] vreg_33_36;
	node n33_36(.left(vreg_32_36), .right(vreg_34_36), .up(vreg_33_37), .down(vreg_33_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_36), .sw(sw));
	wire signed[17:0] vwire_33_37;
	reg signed[17:0] vreg_33_37;
	node n33_37(.left(vreg_32_37), .right(vreg_34_37), .up(vreg_33_38), .down(vreg_33_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_37), .sw(sw));
	wire signed[17:0] vwire_33_38;
	reg signed[17:0] vreg_33_38;
	node n33_38(.left(vreg_32_38), .right(vreg_34_38), .up(vreg_33_39), .down(vreg_33_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_38), .sw(sw));
	wire signed[17:0] vwire_33_39;
	reg signed[17:0] vreg_33_39;
	node n33_39(.left(vreg_32_39), .right(vreg_34_39), .up(vreg_33_40), .down(vreg_33_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_39), .sw(sw));
	wire signed[17:0] vwire_33_40;
	reg signed[17:0] vreg_33_40;
	node n33_40(.left(vreg_32_40), .right(vreg_34_40), .up(vreg_33_41), .down(vreg_33_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_40), .sw(sw));
	wire signed[17:0] vwire_33_41;
	reg signed[17:0] vreg_33_41;
	node n33_41(.left(vreg_32_41), .right(vreg_34_41), .up(vreg_33_42), .down(vreg_33_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_41), .sw(sw));
	wire signed[17:0] vwire_33_42;
	reg signed[17:0] vreg_33_42;
	node n33_42(.left(vreg_32_42), .right(vreg_34_42), .up(vreg_33_43), .down(vreg_33_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_42), .sw(sw));
	wire signed[17:0] vwire_33_43;
	reg signed[17:0] vreg_33_43;
	node n33_43(.left(vreg_32_43), .right(vreg_34_43), .up(vreg_33_44), .down(vreg_33_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_43), .sw(sw));
	wire signed[17:0] vwire_33_44;
	reg signed[17:0] vreg_33_44;
	node n33_44(.left(vreg_32_44), .right(vreg_34_44), .up(vreg_33_45), .down(vreg_33_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_44), .sw(sw));
	wire signed[17:0] vwire_33_45;
	reg signed[17:0] vreg_33_45;
	node n33_45(.left(vreg_32_45), .right(vreg_34_45), .up(vreg_33_46), .down(vreg_33_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_45), .sw(sw));
	wire signed[17:0] vwire_33_46;
	reg signed[17:0] vreg_33_46;
	node n33_46(.left(vreg_32_46), .right(vreg_34_46), .up(vreg_33_47), .down(vreg_33_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_46), .sw(sw));
	wire signed[17:0] vwire_33_47;
	reg signed[17:0] vreg_33_47;
	node n33_47(.left(vreg_32_47), .right(vreg_34_47), .up(vreg_33_48), .down(vreg_33_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_47), .sw(sw));
	wire signed[17:0] vwire_33_48;
	reg signed[17:0] vreg_33_48;
	node n33_48(.left(vreg_32_48), .right(vreg_34_48), .up(vreg_33_49), .down(vreg_33_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_48), .sw(sw));
	wire signed[17:0] vwire_33_49;
	reg signed[17:0] vreg_33_49;
	node n33_49(.left(vreg_32_49), .right(vreg_34_49), .up(18'b0), .down(vreg_33_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_33_49), .sw(sw));
	wire signed[17:0] vwire_34_0;
	reg signed[17:0] vreg_34_0;
	node n34_0(.left(vreg_33_0), .right(vreg_35_0), .up(vreg_34_1), .down(vreg_34_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_0), .sw(sw));
	wire signed[17:0] vwire_34_1;
	reg signed[17:0] vreg_34_1;
	node n34_1(.left(vreg_33_1), .right(vreg_35_1), .up(vreg_34_2), .down(vreg_34_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_1), .sw(sw));
	wire signed[17:0] vwire_34_2;
	reg signed[17:0] vreg_34_2;
	node n34_2(.left(vreg_33_2), .right(vreg_35_2), .up(vreg_34_3), .down(vreg_34_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_2), .sw(sw));
	wire signed[17:0] vwire_34_3;
	reg signed[17:0] vreg_34_3;
	node n34_3(.left(vreg_33_3), .right(vreg_35_3), .up(vreg_34_4), .down(vreg_34_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_3), .sw(sw));
	wire signed[17:0] vwire_34_4;
	reg signed[17:0] vreg_34_4;
	node n34_4(.left(vreg_33_4), .right(vreg_35_4), .up(vreg_34_5), .down(vreg_34_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_4), .sw(sw));
	wire signed[17:0] vwire_34_5;
	reg signed[17:0] vreg_34_5;
	node n34_5(.left(vreg_33_5), .right(vreg_35_5), .up(vreg_34_6), .down(vreg_34_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_5), .sw(sw));
	wire signed[17:0] vwire_34_6;
	reg signed[17:0] vreg_34_6;
	node n34_6(.left(vreg_33_6), .right(vreg_35_6), .up(vreg_34_7), .down(vreg_34_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_6), .sw(sw));
	wire signed[17:0] vwire_34_7;
	reg signed[17:0] vreg_34_7;
	node n34_7(.left(vreg_33_7), .right(vreg_35_7), .up(vreg_34_8), .down(vreg_34_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_7), .sw(sw));
	wire signed[17:0] vwire_34_8;
	reg signed[17:0] vreg_34_8;
	node n34_8(.left(vreg_33_8), .right(vreg_35_8), .up(vreg_34_9), .down(vreg_34_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_8), .sw(sw));
	wire signed[17:0] vwire_34_9;
	reg signed[17:0] vreg_34_9;
	node n34_9(.left(vreg_33_9), .right(vreg_35_9), .up(vreg_34_10), .down(vreg_34_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_9), .sw(sw));
	wire signed[17:0] vwire_34_10;
	reg signed[17:0] vreg_34_10;
	node n34_10(.left(vreg_33_10), .right(vreg_35_10), .up(vreg_34_11), .down(vreg_34_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_10), .sw(sw));
	wire signed[17:0] vwire_34_11;
	reg signed[17:0] vreg_34_11;
	node n34_11(.left(vreg_33_11), .right(vreg_35_11), .up(vreg_34_12), .down(vreg_34_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_11), .sw(sw));
	wire signed[17:0] vwire_34_12;
	reg signed[17:0] vreg_34_12;
	node n34_12(.left(vreg_33_12), .right(vreg_35_12), .up(vreg_34_13), .down(vreg_34_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_12), .sw(sw));
	wire signed[17:0] vwire_34_13;
	reg signed[17:0] vreg_34_13;
	node n34_13(.left(vreg_33_13), .right(vreg_35_13), .up(vreg_34_14), .down(vreg_34_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_13), .sw(sw));
	wire signed[17:0] vwire_34_14;
	reg signed[17:0] vreg_34_14;
	node n34_14(.left(vreg_33_14), .right(vreg_35_14), .up(vreg_34_15), .down(vreg_34_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_14), .sw(sw));
	wire signed[17:0] vwire_34_15;
	reg signed[17:0] vreg_34_15;
	node n34_15(.left(vreg_33_15), .right(vreg_35_15), .up(vreg_34_16), .down(vreg_34_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_15), .sw(sw));
	wire signed[17:0] vwire_34_16;
	reg signed[17:0] vreg_34_16;
	node n34_16(.left(vreg_33_16), .right(vreg_35_16), .up(vreg_34_17), .down(vreg_34_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_16), .sw(sw));
	wire signed[17:0] vwire_34_17;
	reg signed[17:0] vreg_34_17;
	node n34_17(.left(vreg_33_17), .right(vreg_35_17), .up(vreg_34_18), .down(vreg_34_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_17), .sw(sw));
	wire signed[17:0] vwire_34_18;
	reg signed[17:0] vreg_34_18;
	node n34_18(.left(vreg_33_18), .right(vreg_35_18), .up(vreg_34_19), .down(vreg_34_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_18), .sw(sw));
	wire signed[17:0] vwire_34_19;
	reg signed[17:0] vreg_34_19;
	node n34_19(.left(vreg_33_19), .right(vreg_35_19), .up(vreg_34_20), .down(vreg_34_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_19), .sw(sw));
	wire signed[17:0] vwire_34_20;
	reg signed[17:0] vreg_34_20;
	node n34_20(.left(vreg_33_20), .right(vreg_35_20), .up(vreg_34_21), .down(vreg_34_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_20), .sw(sw));
	wire signed[17:0] vwire_34_21;
	reg signed[17:0] vreg_34_21;
	node n34_21(.left(vreg_33_21), .right(vreg_35_21), .up(vreg_34_22), .down(vreg_34_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_21), .sw(sw));
	wire signed[17:0] vwire_34_22;
	reg signed[17:0] vreg_34_22;
	node n34_22(.left(vreg_33_22), .right(vreg_35_22), .up(vreg_34_23), .down(vreg_34_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_22), .sw(sw));
	wire signed[17:0] vwire_34_23;
	reg signed[17:0] vreg_34_23;
	node n34_23(.left(vreg_33_23), .right(vreg_35_23), .up(vreg_34_24), .down(vreg_34_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_23), .sw(sw));
	wire signed[17:0] vwire_34_24;
	reg signed[17:0] vreg_34_24;
	node n34_24(.left(vreg_33_24), .right(vreg_35_24), .up(vreg_34_25), .down(vreg_34_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_24), .sw(sw));
	wire signed[17:0] vwire_34_25;
	reg signed[17:0] vreg_34_25;
	node n34_25(.left(vreg_33_25), .right(vreg_35_25), .up(vreg_34_26), .down(vreg_34_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_25), .sw(sw));
	wire signed[17:0] vwire_34_26;
	reg signed[17:0] vreg_34_26;
	node n34_26(.left(vreg_33_26), .right(vreg_35_26), .up(vreg_34_27), .down(vreg_34_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_26), .sw(sw));
	wire signed[17:0] vwire_34_27;
	reg signed[17:0] vreg_34_27;
	node n34_27(.left(vreg_33_27), .right(vreg_35_27), .up(vreg_34_28), .down(vreg_34_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_27), .sw(sw));
	wire signed[17:0] vwire_34_28;
	reg signed[17:0] vreg_34_28;
	node n34_28(.left(vreg_33_28), .right(vreg_35_28), .up(vreg_34_29), .down(vreg_34_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_28), .sw(sw));
	wire signed[17:0] vwire_34_29;
	reg signed[17:0] vreg_34_29;
	node n34_29(.left(vreg_33_29), .right(vreg_35_29), .up(vreg_34_30), .down(vreg_34_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_29), .sw(sw));
	wire signed[17:0] vwire_34_30;
	reg signed[17:0] vreg_34_30;
	node n34_30(.left(vreg_33_30), .right(vreg_35_30), .up(vreg_34_31), .down(vreg_34_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_30), .sw(sw));
	wire signed[17:0] vwire_34_31;
	reg signed[17:0] vreg_34_31;
	node n34_31(.left(vreg_33_31), .right(vreg_35_31), .up(vreg_34_32), .down(vreg_34_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_31), .sw(sw));
	wire signed[17:0] vwire_34_32;
	reg signed[17:0] vreg_34_32;
	node n34_32(.left(vreg_33_32), .right(vreg_35_32), .up(vreg_34_33), .down(vreg_34_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_32), .sw(sw));
	wire signed[17:0] vwire_34_33;
	reg signed[17:0] vreg_34_33;
	node n34_33(.left(vreg_33_33), .right(vreg_35_33), .up(vreg_34_34), .down(vreg_34_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_33), .sw(sw));
	wire signed[17:0] vwire_34_34;
	reg signed[17:0] vreg_34_34;
	node n34_34(.left(vreg_33_34), .right(vreg_35_34), .up(vreg_34_35), .down(vreg_34_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_34), .sw(sw));
	wire signed[17:0] vwire_34_35;
	reg signed[17:0] vreg_34_35;
	node n34_35(.left(vreg_33_35), .right(vreg_35_35), .up(vreg_34_36), .down(vreg_34_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_35), .sw(sw));
	wire signed[17:0] vwire_34_36;
	reg signed[17:0] vreg_34_36;
	node n34_36(.left(vreg_33_36), .right(vreg_35_36), .up(vreg_34_37), .down(vreg_34_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_36), .sw(sw));
	wire signed[17:0] vwire_34_37;
	reg signed[17:0] vreg_34_37;
	node n34_37(.left(vreg_33_37), .right(vreg_35_37), .up(vreg_34_38), .down(vreg_34_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_37), .sw(sw));
	wire signed[17:0] vwire_34_38;
	reg signed[17:0] vreg_34_38;
	node n34_38(.left(vreg_33_38), .right(vreg_35_38), .up(vreg_34_39), .down(vreg_34_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_38), .sw(sw));
	wire signed[17:0] vwire_34_39;
	reg signed[17:0] vreg_34_39;
	node n34_39(.left(vreg_33_39), .right(vreg_35_39), .up(vreg_34_40), .down(vreg_34_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_39), .sw(sw));
	wire signed[17:0] vwire_34_40;
	reg signed[17:0] vreg_34_40;
	node n34_40(.left(vreg_33_40), .right(vreg_35_40), .up(vreg_34_41), .down(vreg_34_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_40), .sw(sw));
	wire signed[17:0] vwire_34_41;
	reg signed[17:0] vreg_34_41;
	node n34_41(.left(vreg_33_41), .right(vreg_35_41), .up(vreg_34_42), .down(vreg_34_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_41), .sw(sw));
	wire signed[17:0] vwire_34_42;
	reg signed[17:0] vreg_34_42;
	node n34_42(.left(vreg_33_42), .right(vreg_35_42), .up(vreg_34_43), .down(vreg_34_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_42), .sw(sw));
	wire signed[17:0] vwire_34_43;
	reg signed[17:0] vreg_34_43;
	node n34_43(.left(vreg_33_43), .right(vreg_35_43), .up(vreg_34_44), .down(vreg_34_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_43), .sw(sw));
	wire signed[17:0] vwire_34_44;
	reg signed[17:0] vreg_34_44;
	node n34_44(.left(vreg_33_44), .right(vreg_35_44), .up(vreg_34_45), .down(vreg_34_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_44), .sw(sw));
	wire signed[17:0] vwire_34_45;
	reg signed[17:0] vreg_34_45;
	node n34_45(.left(vreg_33_45), .right(vreg_35_45), .up(vreg_34_46), .down(vreg_34_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_45), .sw(sw));
	wire signed[17:0] vwire_34_46;
	reg signed[17:0] vreg_34_46;
	node n34_46(.left(vreg_33_46), .right(vreg_35_46), .up(vreg_34_47), .down(vreg_34_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_46), .sw(sw));
	wire signed[17:0] vwire_34_47;
	reg signed[17:0] vreg_34_47;
	node n34_47(.left(vreg_33_47), .right(vreg_35_47), .up(vreg_34_48), .down(vreg_34_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_47), .sw(sw));
	wire signed[17:0] vwire_34_48;
	reg signed[17:0] vreg_34_48;
	node n34_48(.left(vreg_33_48), .right(vreg_35_48), .up(vreg_34_49), .down(vreg_34_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_48), .sw(sw));
	wire signed[17:0] vwire_34_49;
	reg signed[17:0] vreg_34_49;
	node n34_49(.left(vreg_33_49), .right(vreg_35_49), .up(18'b0), .down(vreg_34_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_34_49), .sw(sw));
	wire signed[17:0] vwire_35_0;
	reg signed[17:0] vreg_35_0;
	node n35_0(.left(vreg_34_0), .right(vreg_36_0), .up(vreg_35_1), .down(vreg_35_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_0), .sw(sw));
	wire signed[17:0] vwire_35_1;
	reg signed[17:0] vreg_35_1;
	node n35_1(.left(vreg_34_1), .right(vreg_36_1), .up(vreg_35_2), .down(vreg_35_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_1), .sw(sw));
	wire signed[17:0] vwire_35_2;
	reg signed[17:0] vreg_35_2;
	node n35_2(.left(vreg_34_2), .right(vreg_36_2), .up(vreg_35_3), .down(vreg_35_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_2), .sw(sw));
	wire signed[17:0] vwire_35_3;
	reg signed[17:0] vreg_35_3;
	node n35_3(.left(vreg_34_3), .right(vreg_36_3), .up(vreg_35_4), .down(vreg_35_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_3), .sw(sw));
	wire signed[17:0] vwire_35_4;
	reg signed[17:0] vreg_35_4;
	node n35_4(.left(vreg_34_4), .right(vreg_36_4), .up(vreg_35_5), .down(vreg_35_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_4), .sw(sw));
	wire signed[17:0] vwire_35_5;
	reg signed[17:0] vreg_35_5;
	node n35_5(.left(vreg_34_5), .right(vreg_36_5), .up(vreg_35_6), .down(vreg_35_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_5), .sw(sw));
	wire signed[17:0] vwire_35_6;
	reg signed[17:0] vreg_35_6;
	node n35_6(.left(vreg_34_6), .right(vreg_36_6), .up(vreg_35_7), .down(vreg_35_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_6), .sw(sw));
	wire signed[17:0] vwire_35_7;
	reg signed[17:0] vreg_35_7;
	node n35_7(.left(vreg_34_7), .right(vreg_36_7), .up(vreg_35_8), .down(vreg_35_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_7), .sw(sw));
	wire signed[17:0] vwire_35_8;
	reg signed[17:0] vreg_35_8;
	node n35_8(.left(vreg_34_8), .right(vreg_36_8), .up(vreg_35_9), .down(vreg_35_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_8), .sw(sw));
	wire signed[17:0] vwire_35_9;
	reg signed[17:0] vreg_35_9;
	node n35_9(.left(vreg_34_9), .right(vreg_36_9), .up(vreg_35_10), .down(vreg_35_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_9), .sw(sw));
	wire signed[17:0] vwire_35_10;
	reg signed[17:0] vreg_35_10;
	node n35_10(.left(vreg_34_10), .right(vreg_36_10), .up(vreg_35_11), .down(vreg_35_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_10), .sw(sw));
	wire signed[17:0] vwire_35_11;
	reg signed[17:0] vreg_35_11;
	node n35_11(.left(vreg_34_11), .right(vreg_36_11), .up(vreg_35_12), .down(vreg_35_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_11), .sw(sw));
	wire signed[17:0] vwire_35_12;
	reg signed[17:0] vreg_35_12;
	node n35_12(.left(vreg_34_12), .right(vreg_36_12), .up(vreg_35_13), .down(vreg_35_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_12), .sw(sw));
	wire signed[17:0] vwire_35_13;
	reg signed[17:0] vreg_35_13;
	node n35_13(.left(vreg_34_13), .right(vreg_36_13), .up(vreg_35_14), .down(vreg_35_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_13), .sw(sw));
	wire signed[17:0] vwire_35_14;
	reg signed[17:0] vreg_35_14;
	node n35_14(.left(vreg_34_14), .right(vreg_36_14), .up(vreg_35_15), .down(vreg_35_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_14), .sw(sw));
	wire signed[17:0] vwire_35_15;
	reg signed[17:0] vreg_35_15;
	node n35_15(.left(vreg_34_15), .right(vreg_36_15), .up(vreg_35_16), .down(vreg_35_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_15), .sw(sw));
	wire signed[17:0] vwire_35_16;
	reg signed[17:0] vreg_35_16;
	node n35_16(.left(vreg_34_16), .right(vreg_36_16), .up(vreg_35_17), .down(vreg_35_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_16), .sw(sw));
	wire signed[17:0] vwire_35_17;
	reg signed[17:0] vreg_35_17;
	node n35_17(.left(vreg_34_17), .right(vreg_36_17), .up(vreg_35_18), .down(vreg_35_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_17), .sw(sw));
	wire signed[17:0] vwire_35_18;
	reg signed[17:0] vreg_35_18;
	node n35_18(.left(vreg_34_18), .right(vreg_36_18), .up(vreg_35_19), .down(vreg_35_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_18), .sw(sw));
	wire signed[17:0] vwire_35_19;
	reg signed[17:0] vreg_35_19;
	node n35_19(.left(vreg_34_19), .right(vreg_36_19), .up(vreg_35_20), .down(vreg_35_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_19), .sw(sw));
	wire signed[17:0] vwire_35_20;
	reg signed[17:0] vreg_35_20;
	node n35_20(.left(vreg_34_20), .right(vreg_36_20), .up(vreg_35_21), .down(vreg_35_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_20), .sw(sw));
	wire signed[17:0] vwire_35_21;
	reg signed[17:0] vreg_35_21;
	node n35_21(.left(vreg_34_21), .right(vreg_36_21), .up(vreg_35_22), .down(vreg_35_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_21), .sw(sw));
	wire signed[17:0] vwire_35_22;
	reg signed[17:0] vreg_35_22;
	node n35_22(.left(vreg_34_22), .right(vreg_36_22), .up(vreg_35_23), .down(vreg_35_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_22), .sw(sw));
	wire signed[17:0] vwire_35_23;
	reg signed[17:0] vreg_35_23;
	node n35_23(.left(vreg_34_23), .right(vreg_36_23), .up(vreg_35_24), .down(vreg_35_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_23), .sw(sw));
	wire signed[17:0] vwire_35_24;
	reg signed[17:0] vreg_35_24;
	node n35_24(.left(vreg_34_24), .right(vreg_36_24), .up(vreg_35_25), .down(vreg_35_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_24), .sw(sw));
	wire signed[17:0] vwire_35_25;
	reg signed[17:0] vreg_35_25;
	node n35_25(.left(vreg_34_25), .right(vreg_36_25), .up(vreg_35_26), .down(vreg_35_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_25), .sw(sw));
	wire signed[17:0] vwire_35_26;
	reg signed[17:0] vreg_35_26;
	node n35_26(.left(vreg_34_26), .right(vreg_36_26), .up(vreg_35_27), .down(vreg_35_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_26), .sw(sw));
	wire signed[17:0] vwire_35_27;
	reg signed[17:0] vreg_35_27;
	node n35_27(.left(vreg_34_27), .right(vreg_36_27), .up(vreg_35_28), .down(vreg_35_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_27), .sw(sw));
	wire signed[17:0] vwire_35_28;
	reg signed[17:0] vreg_35_28;
	node n35_28(.left(vreg_34_28), .right(vreg_36_28), .up(vreg_35_29), .down(vreg_35_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_28), .sw(sw));
	wire signed[17:0] vwire_35_29;
	reg signed[17:0] vreg_35_29;
	node n35_29(.left(vreg_34_29), .right(vreg_36_29), .up(vreg_35_30), .down(vreg_35_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_29), .sw(sw));
	wire signed[17:0] vwire_35_30;
	reg signed[17:0] vreg_35_30;
	node n35_30(.left(vreg_34_30), .right(vreg_36_30), .up(vreg_35_31), .down(vreg_35_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_30), .sw(sw));
	wire signed[17:0] vwire_35_31;
	reg signed[17:0] vreg_35_31;
	node n35_31(.left(vreg_34_31), .right(vreg_36_31), .up(vreg_35_32), .down(vreg_35_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_31), .sw(sw));
	wire signed[17:0] vwire_35_32;
	reg signed[17:0] vreg_35_32;
	node n35_32(.left(vreg_34_32), .right(vreg_36_32), .up(vreg_35_33), .down(vreg_35_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_32), .sw(sw));
	wire signed[17:0] vwire_35_33;
	reg signed[17:0] vreg_35_33;
	node n35_33(.left(vreg_34_33), .right(vreg_36_33), .up(vreg_35_34), .down(vreg_35_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_33), .sw(sw));
	wire signed[17:0] vwire_35_34;
	reg signed[17:0] vreg_35_34;
	node n35_34(.left(vreg_34_34), .right(vreg_36_34), .up(vreg_35_35), .down(vreg_35_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_34), .sw(sw));
	wire signed[17:0] vwire_35_35;
	reg signed[17:0] vreg_35_35;
	node n35_35(.left(vreg_34_35), .right(vreg_36_35), .up(vreg_35_36), .down(vreg_35_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_35), .sw(sw));
	wire signed[17:0] vwire_35_36;
	reg signed[17:0] vreg_35_36;
	node n35_36(.left(vreg_34_36), .right(vreg_36_36), .up(vreg_35_37), .down(vreg_35_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_36), .sw(sw));
	wire signed[17:0] vwire_35_37;
	reg signed[17:0] vreg_35_37;
	node n35_37(.left(vreg_34_37), .right(vreg_36_37), .up(vreg_35_38), .down(vreg_35_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_37), .sw(sw));
	wire signed[17:0] vwire_35_38;
	reg signed[17:0] vreg_35_38;
	node n35_38(.left(vreg_34_38), .right(vreg_36_38), .up(vreg_35_39), .down(vreg_35_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_38), .sw(sw));
	wire signed[17:0] vwire_35_39;
	reg signed[17:0] vreg_35_39;
	node n35_39(.left(vreg_34_39), .right(vreg_36_39), .up(vreg_35_40), .down(vreg_35_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_39), .sw(sw));
	wire signed[17:0] vwire_35_40;
	reg signed[17:0] vreg_35_40;
	node n35_40(.left(vreg_34_40), .right(vreg_36_40), .up(vreg_35_41), .down(vreg_35_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_40), .sw(sw));
	wire signed[17:0] vwire_35_41;
	reg signed[17:0] vreg_35_41;
	node n35_41(.left(vreg_34_41), .right(vreg_36_41), .up(vreg_35_42), .down(vreg_35_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_41), .sw(sw));
	wire signed[17:0] vwire_35_42;
	reg signed[17:0] vreg_35_42;
	node n35_42(.left(vreg_34_42), .right(vreg_36_42), .up(vreg_35_43), .down(vreg_35_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_42), .sw(sw));
	wire signed[17:0] vwire_35_43;
	reg signed[17:0] vreg_35_43;
	node n35_43(.left(vreg_34_43), .right(vreg_36_43), .up(vreg_35_44), .down(vreg_35_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_43), .sw(sw));
	wire signed[17:0] vwire_35_44;
	reg signed[17:0] vreg_35_44;
	node n35_44(.left(vreg_34_44), .right(vreg_36_44), .up(vreg_35_45), .down(vreg_35_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_44), .sw(sw));
	wire signed[17:0] vwire_35_45;
	reg signed[17:0] vreg_35_45;
	node n35_45(.left(vreg_34_45), .right(vreg_36_45), .up(vreg_35_46), .down(vreg_35_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_45), .sw(sw));
	wire signed[17:0] vwire_35_46;
	reg signed[17:0] vreg_35_46;
	node n35_46(.left(vreg_34_46), .right(vreg_36_46), .up(vreg_35_47), .down(vreg_35_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_46), .sw(sw));
	wire signed[17:0] vwire_35_47;
	reg signed[17:0] vreg_35_47;
	node n35_47(.left(vreg_34_47), .right(vreg_36_47), .up(vreg_35_48), .down(vreg_35_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_47), .sw(sw));
	wire signed[17:0] vwire_35_48;
	reg signed[17:0] vreg_35_48;
	node n35_48(.left(vreg_34_48), .right(vreg_36_48), .up(vreg_35_49), .down(vreg_35_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_48), .sw(sw));
	wire signed[17:0] vwire_35_49;
	reg signed[17:0] vreg_35_49;
	node n35_49(.left(vreg_34_49), .right(vreg_36_49), .up(18'b0), .down(vreg_35_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_35_49), .sw(sw));
	wire signed[17:0] vwire_36_0;
	reg signed[17:0] vreg_36_0;
	node n36_0(.left(vreg_35_0), .right(vreg_37_0), .up(vreg_36_1), .down(vreg_36_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_0), .sw(sw));
	wire signed[17:0] vwire_36_1;
	reg signed[17:0] vreg_36_1;
	node n36_1(.left(vreg_35_1), .right(vreg_37_1), .up(vreg_36_2), .down(vreg_36_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_1), .sw(sw));
	wire signed[17:0] vwire_36_2;
	reg signed[17:0] vreg_36_2;
	node n36_2(.left(vreg_35_2), .right(vreg_37_2), .up(vreg_36_3), .down(vreg_36_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_2), .sw(sw));
	wire signed[17:0] vwire_36_3;
	reg signed[17:0] vreg_36_3;
	node n36_3(.left(vreg_35_3), .right(vreg_37_3), .up(vreg_36_4), .down(vreg_36_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_3), .sw(sw));
	wire signed[17:0] vwire_36_4;
	reg signed[17:0] vreg_36_4;
	node n36_4(.left(vreg_35_4), .right(vreg_37_4), .up(vreg_36_5), .down(vreg_36_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_4), .sw(sw));
	wire signed[17:0] vwire_36_5;
	reg signed[17:0] vreg_36_5;
	node n36_5(.left(vreg_35_5), .right(vreg_37_5), .up(vreg_36_6), .down(vreg_36_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_5), .sw(sw));
	wire signed[17:0] vwire_36_6;
	reg signed[17:0] vreg_36_6;
	node n36_6(.left(vreg_35_6), .right(vreg_37_6), .up(vreg_36_7), .down(vreg_36_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_6), .sw(sw));
	wire signed[17:0] vwire_36_7;
	reg signed[17:0] vreg_36_7;
	node n36_7(.left(vreg_35_7), .right(vreg_37_7), .up(vreg_36_8), .down(vreg_36_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_7), .sw(sw));
	wire signed[17:0] vwire_36_8;
	reg signed[17:0] vreg_36_8;
	node n36_8(.left(vreg_35_8), .right(vreg_37_8), .up(vreg_36_9), .down(vreg_36_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_8), .sw(sw));
	wire signed[17:0] vwire_36_9;
	reg signed[17:0] vreg_36_9;
	node n36_9(.left(vreg_35_9), .right(vreg_37_9), .up(vreg_36_10), .down(vreg_36_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_9), .sw(sw));
	wire signed[17:0] vwire_36_10;
	reg signed[17:0] vreg_36_10;
	node n36_10(.left(vreg_35_10), .right(vreg_37_10), .up(vreg_36_11), .down(vreg_36_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_10), .sw(sw));
	wire signed[17:0] vwire_36_11;
	reg signed[17:0] vreg_36_11;
	node n36_11(.left(vreg_35_11), .right(vreg_37_11), .up(vreg_36_12), .down(vreg_36_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_11), .sw(sw));
	wire signed[17:0] vwire_36_12;
	reg signed[17:0] vreg_36_12;
	node n36_12(.left(vreg_35_12), .right(vreg_37_12), .up(vreg_36_13), .down(vreg_36_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_12), .sw(sw));
	wire signed[17:0] vwire_36_13;
	reg signed[17:0] vreg_36_13;
	node n36_13(.left(vreg_35_13), .right(vreg_37_13), .up(vreg_36_14), .down(vreg_36_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_13), .sw(sw));
	wire signed[17:0] vwire_36_14;
	reg signed[17:0] vreg_36_14;
	node n36_14(.left(vreg_35_14), .right(vreg_37_14), .up(vreg_36_15), .down(vreg_36_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_14), .sw(sw));
	wire signed[17:0] vwire_36_15;
	reg signed[17:0] vreg_36_15;
	node n36_15(.left(vreg_35_15), .right(vreg_37_15), .up(vreg_36_16), .down(vreg_36_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_15), .sw(sw));
	wire signed[17:0] vwire_36_16;
	reg signed[17:0] vreg_36_16;
	node n36_16(.left(vreg_35_16), .right(vreg_37_16), .up(vreg_36_17), .down(vreg_36_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_16), .sw(sw));
	wire signed[17:0] vwire_36_17;
	reg signed[17:0] vreg_36_17;
	node n36_17(.left(vreg_35_17), .right(vreg_37_17), .up(vreg_36_18), .down(vreg_36_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_17), .sw(sw));
	wire signed[17:0] vwire_36_18;
	reg signed[17:0] vreg_36_18;
	node n36_18(.left(vreg_35_18), .right(vreg_37_18), .up(vreg_36_19), .down(vreg_36_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_18), .sw(sw));
	wire signed[17:0] vwire_36_19;
	reg signed[17:0] vreg_36_19;
	node n36_19(.left(vreg_35_19), .right(vreg_37_19), .up(vreg_36_20), .down(vreg_36_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_19), .sw(sw));
	wire signed[17:0] vwire_36_20;
	reg signed[17:0] vreg_36_20;
	node n36_20(.left(vreg_35_20), .right(vreg_37_20), .up(vreg_36_21), .down(vreg_36_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_20), .sw(sw));
	wire signed[17:0] vwire_36_21;
	reg signed[17:0] vreg_36_21;
	node n36_21(.left(vreg_35_21), .right(vreg_37_21), .up(vreg_36_22), .down(vreg_36_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_21), .sw(sw));
	wire signed[17:0] vwire_36_22;
	reg signed[17:0] vreg_36_22;
	node n36_22(.left(vreg_35_22), .right(vreg_37_22), .up(vreg_36_23), .down(vreg_36_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_22), .sw(sw));
	wire signed[17:0] vwire_36_23;
	reg signed[17:0] vreg_36_23;
	node n36_23(.left(vreg_35_23), .right(vreg_37_23), .up(vreg_36_24), .down(vreg_36_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_23), .sw(sw));
	wire signed[17:0] vwire_36_24;
	reg signed[17:0] vreg_36_24;
	node n36_24(.left(vreg_35_24), .right(vreg_37_24), .up(vreg_36_25), .down(vreg_36_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_24), .sw(sw));
	wire signed[17:0] vwire_36_25;
	reg signed[17:0] vreg_36_25;
	node n36_25(.left(vreg_35_25), .right(vreg_37_25), .up(vreg_36_26), .down(vreg_36_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_25), .sw(sw));
	wire signed[17:0] vwire_36_26;
	reg signed[17:0] vreg_36_26;
	node n36_26(.left(vreg_35_26), .right(vreg_37_26), .up(vreg_36_27), .down(vreg_36_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_26), .sw(sw));
	wire signed[17:0] vwire_36_27;
	reg signed[17:0] vreg_36_27;
	node n36_27(.left(vreg_35_27), .right(vreg_37_27), .up(vreg_36_28), .down(vreg_36_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_27), .sw(sw));
	wire signed[17:0] vwire_36_28;
	reg signed[17:0] vreg_36_28;
	node n36_28(.left(vreg_35_28), .right(vreg_37_28), .up(vreg_36_29), .down(vreg_36_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_28), .sw(sw));
	wire signed[17:0] vwire_36_29;
	reg signed[17:0] vreg_36_29;
	node n36_29(.left(vreg_35_29), .right(vreg_37_29), .up(vreg_36_30), .down(vreg_36_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_29), .sw(sw));
	wire signed[17:0] vwire_36_30;
	reg signed[17:0] vreg_36_30;
	node n36_30(.left(vreg_35_30), .right(vreg_37_30), .up(vreg_36_31), .down(vreg_36_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_30), .sw(sw));
	wire signed[17:0] vwire_36_31;
	reg signed[17:0] vreg_36_31;
	node n36_31(.left(vreg_35_31), .right(vreg_37_31), .up(vreg_36_32), .down(vreg_36_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_31), .sw(sw));
	wire signed[17:0] vwire_36_32;
	reg signed[17:0] vreg_36_32;
	node n36_32(.left(vreg_35_32), .right(vreg_37_32), .up(vreg_36_33), .down(vreg_36_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_32), .sw(sw));
	wire signed[17:0] vwire_36_33;
	reg signed[17:0] vreg_36_33;
	node n36_33(.left(vreg_35_33), .right(vreg_37_33), .up(vreg_36_34), .down(vreg_36_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_33), .sw(sw));
	wire signed[17:0] vwire_36_34;
	reg signed[17:0] vreg_36_34;
	node n36_34(.left(vreg_35_34), .right(vreg_37_34), .up(vreg_36_35), .down(vreg_36_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_34), .sw(sw));
	wire signed[17:0] vwire_36_35;
	reg signed[17:0] vreg_36_35;
	node n36_35(.left(vreg_35_35), .right(vreg_37_35), .up(vreg_36_36), .down(vreg_36_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_35), .sw(sw));
	wire signed[17:0] vwire_36_36;
	reg signed[17:0] vreg_36_36;
	node n36_36(.left(vreg_35_36), .right(vreg_37_36), .up(vreg_36_37), .down(vreg_36_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_36), .sw(sw));
	wire signed[17:0] vwire_36_37;
	reg signed[17:0] vreg_36_37;
	node n36_37(.left(vreg_35_37), .right(vreg_37_37), .up(vreg_36_38), .down(vreg_36_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_37), .sw(sw));
	wire signed[17:0] vwire_36_38;
	reg signed[17:0] vreg_36_38;
	node n36_38(.left(vreg_35_38), .right(vreg_37_38), .up(vreg_36_39), .down(vreg_36_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_38), .sw(sw));
	wire signed[17:0] vwire_36_39;
	reg signed[17:0] vreg_36_39;
	node n36_39(.left(vreg_35_39), .right(vreg_37_39), .up(vreg_36_40), .down(vreg_36_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_39), .sw(sw));
	wire signed[17:0] vwire_36_40;
	reg signed[17:0] vreg_36_40;
	node n36_40(.left(vreg_35_40), .right(vreg_37_40), .up(vreg_36_41), .down(vreg_36_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_40), .sw(sw));
	wire signed[17:0] vwire_36_41;
	reg signed[17:0] vreg_36_41;
	node n36_41(.left(vreg_35_41), .right(vreg_37_41), .up(vreg_36_42), .down(vreg_36_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_41), .sw(sw));
	wire signed[17:0] vwire_36_42;
	reg signed[17:0] vreg_36_42;
	node n36_42(.left(vreg_35_42), .right(vreg_37_42), .up(vreg_36_43), .down(vreg_36_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_42), .sw(sw));
	wire signed[17:0] vwire_36_43;
	reg signed[17:0] vreg_36_43;
	node n36_43(.left(vreg_35_43), .right(vreg_37_43), .up(vreg_36_44), .down(vreg_36_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_43), .sw(sw));
	wire signed[17:0] vwire_36_44;
	reg signed[17:0] vreg_36_44;
	node n36_44(.left(vreg_35_44), .right(vreg_37_44), .up(vreg_36_45), .down(vreg_36_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_44), .sw(sw));
	wire signed[17:0] vwire_36_45;
	reg signed[17:0] vreg_36_45;
	node n36_45(.left(vreg_35_45), .right(vreg_37_45), .up(vreg_36_46), .down(vreg_36_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_45), .sw(sw));
	wire signed[17:0] vwire_36_46;
	reg signed[17:0] vreg_36_46;
	node n36_46(.left(vreg_35_46), .right(vreg_37_46), .up(vreg_36_47), .down(vreg_36_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_46), .sw(sw));
	wire signed[17:0] vwire_36_47;
	reg signed[17:0] vreg_36_47;
	node n36_47(.left(vreg_35_47), .right(vreg_37_47), .up(vreg_36_48), .down(vreg_36_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_47), .sw(sw));
	wire signed[17:0] vwire_36_48;
	reg signed[17:0] vreg_36_48;
	node n36_48(.left(vreg_35_48), .right(vreg_37_48), .up(vreg_36_49), .down(vreg_36_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_48), .sw(sw));
	wire signed[17:0] vwire_36_49;
	reg signed[17:0] vreg_36_49;
	node n36_49(.left(vreg_35_49), .right(vreg_37_49), .up(18'b0), .down(vreg_36_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_36_49), .sw(sw));
	wire signed[17:0] vwire_37_0;
	reg signed[17:0] vreg_37_0;
	node n37_0(.left(vreg_36_0), .right(vreg_38_0), .up(vreg_37_1), .down(vreg_37_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_0), .sw(sw));
	wire signed[17:0] vwire_37_1;
	reg signed[17:0] vreg_37_1;
	node n37_1(.left(vreg_36_1), .right(vreg_38_1), .up(vreg_37_2), .down(vreg_37_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_1), .sw(sw));
	wire signed[17:0] vwire_37_2;
	reg signed[17:0] vreg_37_2;
	node n37_2(.left(vreg_36_2), .right(vreg_38_2), .up(vreg_37_3), .down(vreg_37_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_2), .sw(sw));
	wire signed[17:0] vwire_37_3;
	reg signed[17:0] vreg_37_3;
	node n37_3(.left(vreg_36_3), .right(vreg_38_3), .up(vreg_37_4), .down(vreg_37_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_3), .sw(sw));
	wire signed[17:0] vwire_37_4;
	reg signed[17:0] vreg_37_4;
	node n37_4(.left(vreg_36_4), .right(vreg_38_4), .up(vreg_37_5), .down(vreg_37_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_4), .sw(sw));
	wire signed[17:0] vwire_37_5;
	reg signed[17:0] vreg_37_5;
	node n37_5(.left(vreg_36_5), .right(vreg_38_5), .up(vreg_37_6), .down(vreg_37_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_5), .sw(sw));
	wire signed[17:0] vwire_37_6;
	reg signed[17:0] vreg_37_6;
	node n37_6(.left(vreg_36_6), .right(vreg_38_6), .up(vreg_37_7), .down(vreg_37_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_6), .sw(sw));
	wire signed[17:0] vwire_37_7;
	reg signed[17:0] vreg_37_7;
	node n37_7(.left(vreg_36_7), .right(vreg_38_7), .up(vreg_37_8), .down(vreg_37_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_7), .sw(sw));
	wire signed[17:0] vwire_37_8;
	reg signed[17:0] vreg_37_8;
	node n37_8(.left(vreg_36_8), .right(vreg_38_8), .up(vreg_37_9), .down(vreg_37_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_8), .sw(sw));
	wire signed[17:0] vwire_37_9;
	reg signed[17:0] vreg_37_9;
	node n37_9(.left(vreg_36_9), .right(vreg_38_9), .up(vreg_37_10), .down(vreg_37_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_9), .sw(sw));
	wire signed[17:0] vwire_37_10;
	reg signed[17:0] vreg_37_10;
	node n37_10(.left(vreg_36_10), .right(vreg_38_10), .up(vreg_37_11), .down(vreg_37_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_10), .sw(sw));
	wire signed[17:0] vwire_37_11;
	reg signed[17:0] vreg_37_11;
	node n37_11(.left(vreg_36_11), .right(vreg_38_11), .up(vreg_37_12), .down(vreg_37_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_11), .sw(sw));
	wire signed[17:0] vwire_37_12;
	reg signed[17:0] vreg_37_12;
	node n37_12(.left(vreg_36_12), .right(vreg_38_12), .up(vreg_37_13), .down(vreg_37_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_12), .sw(sw));
	wire signed[17:0] vwire_37_13;
	reg signed[17:0] vreg_37_13;
	node n37_13(.left(vreg_36_13), .right(vreg_38_13), .up(vreg_37_14), .down(vreg_37_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_13), .sw(sw));
	wire signed[17:0] vwire_37_14;
	reg signed[17:0] vreg_37_14;
	node n37_14(.left(vreg_36_14), .right(vreg_38_14), .up(vreg_37_15), .down(vreg_37_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_14), .sw(sw));
	wire signed[17:0] vwire_37_15;
	reg signed[17:0] vreg_37_15;
	node n37_15(.left(vreg_36_15), .right(vreg_38_15), .up(vreg_37_16), .down(vreg_37_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_15), .sw(sw));
	wire signed[17:0] vwire_37_16;
	reg signed[17:0] vreg_37_16;
	node n37_16(.left(vreg_36_16), .right(vreg_38_16), .up(vreg_37_17), .down(vreg_37_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_16), .sw(sw));
	wire signed[17:0] vwire_37_17;
	reg signed[17:0] vreg_37_17;
	node n37_17(.left(vreg_36_17), .right(vreg_38_17), .up(vreg_37_18), .down(vreg_37_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_17), .sw(sw));
	wire signed[17:0] vwire_37_18;
	reg signed[17:0] vreg_37_18;
	node n37_18(.left(vreg_36_18), .right(vreg_38_18), .up(vreg_37_19), .down(vreg_37_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_18), .sw(sw));
	wire signed[17:0] vwire_37_19;
	reg signed[17:0] vreg_37_19;
	node n37_19(.left(vreg_36_19), .right(vreg_38_19), .up(vreg_37_20), .down(vreg_37_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_19), .sw(sw));
	wire signed[17:0] vwire_37_20;
	reg signed[17:0] vreg_37_20;
	node n37_20(.left(vreg_36_20), .right(vreg_38_20), .up(vreg_37_21), .down(vreg_37_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_20), .sw(sw));
	wire signed[17:0] vwire_37_21;
	reg signed[17:0] vreg_37_21;
	node n37_21(.left(vreg_36_21), .right(vreg_38_21), .up(vreg_37_22), .down(vreg_37_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_21), .sw(sw));
	wire signed[17:0] vwire_37_22;
	reg signed[17:0] vreg_37_22;
	node n37_22(.left(vreg_36_22), .right(vreg_38_22), .up(vreg_37_23), .down(vreg_37_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_22), .sw(sw));
	wire signed[17:0] vwire_37_23;
	reg signed[17:0] vreg_37_23;
	node n37_23(.left(vreg_36_23), .right(vreg_38_23), .up(vreg_37_24), .down(vreg_37_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_23), .sw(sw));
	wire signed[17:0] vwire_37_24;
	reg signed[17:0] vreg_37_24;
	node n37_24(.left(vreg_36_24), .right(vreg_38_24), .up(vreg_37_25), .down(vreg_37_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_24), .sw(sw));
	wire signed[17:0] vwire_37_25;
	reg signed[17:0] vreg_37_25;
	node n37_25(.left(vreg_36_25), .right(vreg_38_25), .up(vreg_37_26), .down(vreg_37_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_25), .sw(sw));
	wire signed[17:0] vwire_37_26;
	reg signed[17:0] vreg_37_26;
	node n37_26(.left(vreg_36_26), .right(vreg_38_26), .up(vreg_37_27), .down(vreg_37_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_26), .sw(sw));
	wire signed[17:0] vwire_37_27;
	reg signed[17:0] vreg_37_27;
	node n37_27(.left(vreg_36_27), .right(vreg_38_27), .up(vreg_37_28), .down(vreg_37_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_27), .sw(sw));
	wire signed[17:0] vwire_37_28;
	reg signed[17:0] vreg_37_28;
	node n37_28(.left(vreg_36_28), .right(vreg_38_28), .up(vreg_37_29), .down(vreg_37_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_28), .sw(sw));
	wire signed[17:0] vwire_37_29;
	reg signed[17:0] vreg_37_29;
	node n37_29(.left(vreg_36_29), .right(vreg_38_29), .up(vreg_37_30), .down(vreg_37_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_29), .sw(sw));
	wire signed[17:0] vwire_37_30;
	reg signed[17:0] vreg_37_30;
	node n37_30(.left(vreg_36_30), .right(vreg_38_30), .up(vreg_37_31), .down(vreg_37_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_30), .sw(sw));
	wire signed[17:0] vwire_37_31;
	reg signed[17:0] vreg_37_31;
	node n37_31(.left(vreg_36_31), .right(vreg_38_31), .up(vreg_37_32), .down(vreg_37_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_31), .sw(sw));
	wire signed[17:0] vwire_37_32;
	reg signed[17:0] vreg_37_32;
	node n37_32(.left(vreg_36_32), .right(vreg_38_32), .up(vreg_37_33), .down(vreg_37_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_32), .sw(sw));
	wire signed[17:0] vwire_37_33;
	reg signed[17:0] vreg_37_33;
	node n37_33(.left(vreg_36_33), .right(vreg_38_33), .up(vreg_37_34), .down(vreg_37_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_33), .sw(sw));
	wire signed[17:0] vwire_37_34;
	reg signed[17:0] vreg_37_34;
	node n37_34(.left(vreg_36_34), .right(vreg_38_34), .up(vreg_37_35), .down(vreg_37_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_34), .sw(sw));
	wire signed[17:0] vwire_37_35;
	reg signed[17:0] vreg_37_35;
	node n37_35(.left(vreg_36_35), .right(vreg_38_35), .up(vreg_37_36), .down(vreg_37_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_35), .sw(sw));
	wire signed[17:0] vwire_37_36;
	reg signed[17:0] vreg_37_36;
	node n37_36(.left(vreg_36_36), .right(vreg_38_36), .up(vreg_37_37), .down(vreg_37_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_36), .sw(sw));
	wire signed[17:0] vwire_37_37;
	reg signed[17:0] vreg_37_37;
	node n37_37(.left(vreg_36_37), .right(vreg_38_37), .up(vreg_37_38), .down(vreg_37_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_37), .sw(sw));
	wire signed[17:0] vwire_37_38;
	reg signed[17:0] vreg_37_38;
	node n37_38(.left(vreg_36_38), .right(vreg_38_38), .up(vreg_37_39), .down(vreg_37_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_38), .sw(sw));
	wire signed[17:0] vwire_37_39;
	reg signed[17:0] vreg_37_39;
	node n37_39(.left(vreg_36_39), .right(vreg_38_39), .up(vreg_37_40), .down(vreg_37_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_39), .sw(sw));
	wire signed[17:0] vwire_37_40;
	reg signed[17:0] vreg_37_40;
	node n37_40(.left(vreg_36_40), .right(vreg_38_40), .up(vreg_37_41), .down(vreg_37_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_40), .sw(sw));
	wire signed[17:0] vwire_37_41;
	reg signed[17:0] vreg_37_41;
	node n37_41(.left(vreg_36_41), .right(vreg_38_41), .up(vreg_37_42), .down(vreg_37_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_41), .sw(sw));
	wire signed[17:0] vwire_37_42;
	reg signed[17:0] vreg_37_42;
	node n37_42(.left(vreg_36_42), .right(vreg_38_42), .up(vreg_37_43), .down(vreg_37_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_42), .sw(sw));
	wire signed[17:0] vwire_37_43;
	reg signed[17:0] vreg_37_43;
	node n37_43(.left(vreg_36_43), .right(vreg_38_43), .up(vreg_37_44), .down(vreg_37_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_43), .sw(sw));
	wire signed[17:0] vwire_37_44;
	reg signed[17:0] vreg_37_44;
	node n37_44(.left(vreg_36_44), .right(vreg_38_44), .up(vreg_37_45), .down(vreg_37_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_44), .sw(sw));
	wire signed[17:0] vwire_37_45;
	reg signed[17:0] vreg_37_45;
	node n37_45(.left(vreg_36_45), .right(vreg_38_45), .up(vreg_37_46), .down(vreg_37_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_45), .sw(sw));
	wire signed[17:0] vwire_37_46;
	reg signed[17:0] vreg_37_46;
	node n37_46(.left(vreg_36_46), .right(vreg_38_46), .up(vreg_37_47), .down(vreg_37_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_46), .sw(sw));
	wire signed[17:0] vwire_37_47;
	reg signed[17:0] vreg_37_47;
	node n37_47(.left(vreg_36_47), .right(vreg_38_47), .up(vreg_37_48), .down(vreg_37_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_47), .sw(sw));
	wire signed[17:0] vwire_37_48;
	reg signed[17:0] vreg_37_48;
	node n37_48(.left(vreg_36_48), .right(vreg_38_48), .up(vreg_37_49), .down(vreg_37_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_48), .sw(sw));
	wire signed[17:0] vwire_37_49;
	reg signed[17:0] vreg_37_49;
	node n37_49(.left(vreg_36_49), .right(vreg_38_49), .up(18'b0), .down(vreg_37_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_37_49), .sw(sw));
	wire signed[17:0] vwire_38_0;
	reg signed[17:0] vreg_38_0;
	node n38_0(.left(vreg_37_0), .right(vreg_39_0), .up(vreg_38_1), .down(vreg_38_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_0), .sw(sw));
	wire signed[17:0] vwire_38_1;
	reg signed[17:0] vreg_38_1;
	node n38_1(.left(vreg_37_1), .right(vreg_39_1), .up(vreg_38_2), .down(vreg_38_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_1), .sw(sw));
	wire signed[17:0] vwire_38_2;
	reg signed[17:0] vreg_38_2;
	node n38_2(.left(vreg_37_2), .right(vreg_39_2), .up(vreg_38_3), .down(vreg_38_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_2), .sw(sw));
	wire signed[17:0] vwire_38_3;
	reg signed[17:0] vreg_38_3;
	node n38_3(.left(vreg_37_3), .right(vreg_39_3), .up(vreg_38_4), .down(vreg_38_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_3), .sw(sw));
	wire signed[17:0] vwire_38_4;
	reg signed[17:0] vreg_38_4;
	node n38_4(.left(vreg_37_4), .right(vreg_39_4), .up(vreg_38_5), .down(vreg_38_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_4), .sw(sw));
	wire signed[17:0] vwire_38_5;
	reg signed[17:0] vreg_38_5;
	node n38_5(.left(vreg_37_5), .right(vreg_39_5), .up(vreg_38_6), .down(vreg_38_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_5), .sw(sw));
	wire signed[17:0] vwire_38_6;
	reg signed[17:0] vreg_38_6;
	node n38_6(.left(vreg_37_6), .right(vreg_39_6), .up(vreg_38_7), .down(vreg_38_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_6), .sw(sw));
	wire signed[17:0] vwire_38_7;
	reg signed[17:0] vreg_38_7;
	node n38_7(.left(vreg_37_7), .right(vreg_39_7), .up(vreg_38_8), .down(vreg_38_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_7), .sw(sw));
	wire signed[17:0] vwire_38_8;
	reg signed[17:0] vreg_38_8;
	node n38_8(.left(vreg_37_8), .right(vreg_39_8), .up(vreg_38_9), .down(vreg_38_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_8), .sw(sw));
	wire signed[17:0] vwire_38_9;
	reg signed[17:0] vreg_38_9;
	node n38_9(.left(vreg_37_9), .right(vreg_39_9), .up(vreg_38_10), .down(vreg_38_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_9), .sw(sw));
	wire signed[17:0] vwire_38_10;
	reg signed[17:0] vreg_38_10;
	node n38_10(.left(vreg_37_10), .right(vreg_39_10), .up(vreg_38_11), .down(vreg_38_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_10), .sw(sw));
	wire signed[17:0] vwire_38_11;
	reg signed[17:0] vreg_38_11;
	node n38_11(.left(vreg_37_11), .right(vreg_39_11), .up(vreg_38_12), .down(vreg_38_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_11), .sw(sw));
	wire signed[17:0] vwire_38_12;
	reg signed[17:0] vreg_38_12;
	node n38_12(.left(vreg_37_12), .right(vreg_39_12), .up(vreg_38_13), .down(vreg_38_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_12), .sw(sw));
	wire signed[17:0] vwire_38_13;
	reg signed[17:0] vreg_38_13;
	node n38_13(.left(vreg_37_13), .right(vreg_39_13), .up(vreg_38_14), .down(vreg_38_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_13), .sw(sw));
	wire signed[17:0] vwire_38_14;
	reg signed[17:0] vreg_38_14;
	node n38_14(.left(vreg_37_14), .right(vreg_39_14), .up(vreg_38_15), .down(vreg_38_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_14), .sw(sw));
	wire signed[17:0] vwire_38_15;
	reg signed[17:0] vreg_38_15;
	node n38_15(.left(vreg_37_15), .right(vreg_39_15), .up(vreg_38_16), .down(vreg_38_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_15), .sw(sw));
	wire signed[17:0] vwire_38_16;
	reg signed[17:0] vreg_38_16;
	node n38_16(.left(vreg_37_16), .right(vreg_39_16), .up(vreg_38_17), .down(vreg_38_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_16), .sw(sw));
	wire signed[17:0] vwire_38_17;
	reg signed[17:0] vreg_38_17;
	node n38_17(.left(vreg_37_17), .right(vreg_39_17), .up(vreg_38_18), .down(vreg_38_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_17), .sw(sw));
	wire signed[17:0] vwire_38_18;
	reg signed[17:0] vreg_38_18;
	node n38_18(.left(vreg_37_18), .right(vreg_39_18), .up(vreg_38_19), .down(vreg_38_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_18), .sw(sw));
	wire signed[17:0] vwire_38_19;
	reg signed[17:0] vreg_38_19;
	node n38_19(.left(vreg_37_19), .right(vreg_39_19), .up(vreg_38_20), .down(vreg_38_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_19), .sw(sw));
	wire signed[17:0] vwire_38_20;
	reg signed[17:0] vreg_38_20;
	node n38_20(.left(vreg_37_20), .right(vreg_39_20), .up(vreg_38_21), .down(vreg_38_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_20), .sw(sw));
	wire signed[17:0] vwire_38_21;
	reg signed[17:0] vreg_38_21;
	node n38_21(.left(vreg_37_21), .right(vreg_39_21), .up(vreg_38_22), .down(vreg_38_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_21), .sw(sw));
	wire signed[17:0] vwire_38_22;
	reg signed[17:0] vreg_38_22;
	node n38_22(.left(vreg_37_22), .right(vreg_39_22), .up(vreg_38_23), .down(vreg_38_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_22), .sw(sw));
	wire signed[17:0] vwire_38_23;
	reg signed[17:0] vreg_38_23;
	node n38_23(.left(vreg_37_23), .right(vreg_39_23), .up(vreg_38_24), .down(vreg_38_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_23), .sw(sw));
	wire signed[17:0] vwire_38_24;
	reg signed[17:0] vreg_38_24;
	node n38_24(.left(vreg_37_24), .right(vreg_39_24), .up(vreg_38_25), .down(vreg_38_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_24), .sw(sw));
	wire signed[17:0] vwire_38_25;
	reg signed[17:0] vreg_38_25;
	node n38_25(.left(vreg_37_25), .right(vreg_39_25), .up(vreg_38_26), .down(vreg_38_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_25), .sw(sw));
	wire signed[17:0] vwire_38_26;
	reg signed[17:0] vreg_38_26;
	node n38_26(.left(vreg_37_26), .right(vreg_39_26), .up(vreg_38_27), .down(vreg_38_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_26), .sw(sw));
	wire signed[17:0] vwire_38_27;
	reg signed[17:0] vreg_38_27;
	node n38_27(.left(vreg_37_27), .right(vreg_39_27), .up(vreg_38_28), .down(vreg_38_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_27), .sw(sw));
	wire signed[17:0] vwire_38_28;
	reg signed[17:0] vreg_38_28;
	node n38_28(.left(vreg_37_28), .right(vreg_39_28), .up(vreg_38_29), .down(vreg_38_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_28), .sw(sw));
	wire signed[17:0] vwire_38_29;
	reg signed[17:0] vreg_38_29;
	node n38_29(.left(vreg_37_29), .right(vreg_39_29), .up(vreg_38_30), .down(vreg_38_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_29), .sw(sw));
	wire signed[17:0] vwire_38_30;
	reg signed[17:0] vreg_38_30;
	node n38_30(.left(vreg_37_30), .right(vreg_39_30), .up(vreg_38_31), .down(vreg_38_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_30), .sw(sw));
	wire signed[17:0] vwire_38_31;
	reg signed[17:0] vreg_38_31;
	node n38_31(.left(vreg_37_31), .right(vreg_39_31), .up(vreg_38_32), .down(vreg_38_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_31), .sw(sw));
	wire signed[17:0] vwire_38_32;
	reg signed[17:0] vreg_38_32;
	node n38_32(.left(vreg_37_32), .right(vreg_39_32), .up(vreg_38_33), .down(vreg_38_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_32), .sw(sw));
	wire signed[17:0] vwire_38_33;
	reg signed[17:0] vreg_38_33;
	node n38_33(.left(vreg_37_33), .right(vreg_39_33), .up(vreg_38_34), .down(vreg_38_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_33), .sw(sw));
	wire signed[17:0] vwire_38_34;
	reg signed[17:0] vreg_38_34;
	node n38_34(.left(vreg_37_34), .right(vreg_39_34), .up(vreg_38_35), .down(vreg_38_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_34), .sw(sw));
	wire signed[17:0] vwire_38_35;
	reg signed[17:0] vreg_38_35;
	node n38_35(.left(vreg_37_35), .right(vreg_39_35), .up(vreg_38_36), .down(vreg_38_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_35), .sw(sw));
	wire signed[17:0] vwire_38_36;
	reg signed[17:0] vreg_38_36;
	node n38_36(.left(vreg_37_36), .right(vreg_39_36), .up(vreg_38_37), .down(vreg_38_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_36), .sw(sw));
	wire signed[17:0] vwire_38_37;
	reg signed[17:0] vreg_38_37;
	node n38_37(.left(vreg_37_37), .right(vreg_39_37), .up(vreg_38_38), .down(vreg_38_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_37), .sw(sw));
	wire signed[17:0] vwire_38_38;
	reg signed[17:0] vreg_38_38;
	node n38_38(.left(vreg_37_38), .right(vreg_39_38), .up(vreg_38_39), .down(vreg_38_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_38), .sw(sw));
	wire signed[17:0] vwire_38_39;
	reg signed[17:0] vreg_38_39;
	node n38_39(.left(vreg_37_39), .right(vreg_39_39), .up(vreg_38_40), .down(vreg_38_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_39), .sw(sw));
	wire signed[17:0] vwire_38_40;
	reg signed[17:0] vreg_38_40;
	node n38_40(.left(vreg_37_40), .right(vreg_39_40), .up(vreg_38_41), .down(vreg_38_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_40), .sw(sw));
	wire signed[17:0] vwire_38_41;
	reg signed[17:0] vreg_38_41;
	node n38_41(.left(vreg_37_41), .right(vreg_39_41), .up(vreg_38_42), .down(vreg_38_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_41), .sw(sw));
	wire signed[17:0] vwire_38_42;
	reg signed[17:0] vreg_38_42;
	node n38_42(.left(vreg_37_42), .right(vreg_39_42), .up(vreg_38_43), .down(vreg_38_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_42), .sw(sw));
	wire signed[17:0] vwire_38_43;
	reg signed[17:0] vreg_38_43;
	node n38_43(.left(vreg_37_43), .right(vreg_39_43), .up(vreg_38_44), .down(vreg_38_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_43), .sw(sw));
	wire signed[17:0] vwire_38_44;
	reg signed[17:0] vreg_38_44;
	node n38_44(.left(vreg_37_44), .right(vreg_39_44), .up(vreg_38_45), .down(vreg_38_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_44), .sw(sw));
	wire signed[17:0] vwire_38_45;
	reg signed[17:0] vreg_38_45;
	node n38_45(.left(vreg_37_45), .right(vreg_39_45), .up(vreg_38_46), .down(vreg_38_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_45), .sw(sw));
	wire signed[17:0] vwire_38_46;
	reg signed[17:0] vreg_38_46;
	node n38_46(.left(vreg_37_46), .right(vreg_39_46), .up(vreg_38_47), .down(vreg_38_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_46), .sw(sw));
	wire signed[17:0] vwire_38_47;
	reg signed[17:0] vreg_38_47;
	node n38_47(.left(vreg_37_47), .right(vreg_39_47), .up(vreg_38_48), .down(vreg_38_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_47), .sw(sw));
	wire signed[17:0] vwire_38_48;
	reg signed[17:0] vreg_38_48;
	node n38_48(.left(vreg_37_48), .right(vreg_39_48), .up(vreg_38_49), .down(vreg_38_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_48), .sw(sw));
	wire signed[17:0] vwire_38_49;
	reg signed[17:0] vreg_38_49;
	node n38_49(.left(vreg_37_49), .right(vreg_39_49), .up(18'b0), .down(vreg_38_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_38_49), .sw(sw));
	wire signed[17:0] vwire_39_0;
	reg signed[17:0] vreg_39_0;
	node n39_0(.left(vreg_38_0), .right(vreg_40_0), .up(vreg_39_1), .down(vreg_39_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_0), .sw(sw));
	wire signed[17:0] vwire_39_1;
	reg signed[17:0] vreg_39_1;
	node n39_1(.left(vreg_38_1), .right(vreg_40_1), .up(vreg_39_2), .down(vreg_39_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_1), .sw(sw));
	wire signed[17:0] vwire_39_2;
	reg signed[17:0] vreg_39_2;
	node n39_2(.left(vreg_38_2), .right(vreg_40_2), .up(vreg_39_3), .down(vreg_39_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_2), .sw(sw));
	wire signed[17:0] vwire_39_3;
	reg signed[17:0] vreg_39_3;
	node n39_3(.left(vreg_38_3), .right(vreg_40_3), .up(vreg_39_4), .down(vreg_39_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_3), .sw(sw));
	wire signed[17:0] vwire_39_4;
	reg signed[17:0] vreg_39_4;
	node n39_4(.left(vreg_38_4), .right(vreg_40_4), .up(vreg_39_5), .down(vreg_39_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_4), .sw(sw));
	wire signed[17:0] vwire_39_5;
	reg signed[17:0] vreg_39_5;
	node n39_5(.left(vreg_38_5), .right(vreg_40_5), .up(vreg_39_6), .down(vreg_39_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_5), .sw(sw));
	wire signed[17:0] vwire_39_6;
	reg signed[17:0] vreg_39_6;
	node n39_6(.left(vreg_38_6), .right(vreg_40_6), .up(vreg_39_7), .down(vreg_39_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_6), .sw(sw));
	wire signed[17:0] vwire_39_7;
	reg signed[17:0] vreg_39_7;
	node n39_7(.left(vreg_38_7), .right(vreg_40_7), .up(vreg_39_8), .down(vreg_39_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_7), .sw(sw));
	wire signed[17:0] vwire_39_8;
	reg signed[17:0] vreg_39_8;
	node n39_8(.left(vreg_38_8), .right(vreg_40_8), .up(vreg_39_9), .down(vreg_39_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_8), .sw(sw));
	wire signed[17:0] vwire_39_9;
	reg signed[17:0] vreg_39_9;
	node n39_9(.left(vreg_38_9), .right(vreg_40_9), .up(vreg_39_10), .down(vreg_39_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_9), .sw(sw));
	wire signed[17:0] vwire_39_10;
	reg signed[17:0] vreg_39_10;
	node n39_10(.left(vreg_38_10), .right(vreg_40_10), .up(vreg_39_11), .down(vreg_39_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_10), .sw(sw));
	wire signed[17:0] vwire_39_11;
	reg signed[17:0] vreg_39_11;
	node n39_11(.left(vreg_38_11), .right(vreg_40_11), .up(vreg_39_12), .down(vreg_39_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_11), .sw(sw));
	wire signed[17:0] vwire_39_12;
	reg signed[17:0] vreg_39_12;
	node n39_12(.left(vreg_38_12), .right(vreg_40_12), .up(vreg_39_13), .down(vreg_39_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_12), .sw(sw));
	wire signed[17:0] vwire_39_13;
	reg signed[17:0] vreg_39_13;
	node n39_13(.left(vreg_38_13), .right(vreg_40_13), .up(vreg_39_14), .down(vreg_39_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_13), .sw(sw));
	wire signed[17:0] vwire_39_14;
	reg signed[17:0] vreg_39_14;
	node n39_14(.left(vreg_38_14), .right(vreg_40_14), .up(vreg_39_15), .down(vreg_39_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_14), .sw(sw));
	wire signed[17:0] vwire_39_15;
	reg signed[17:0] vreg_39_15;
	node n39_15(.left(vreg_38_15), .right(vreg_40_15), .up(vreg_39_16), .down(vreg_39_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_15), .sw(sw));
	wire signed[17:0] vwire_39_16;
	reg signed[17:0] vreg_39_16;
	node n39_16(.left(vreg_38_16), .right(vreg_40_16), .up(vreg_39_17), .down(vreg_39_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_16), .sw(sw));
	wire signed[17:0] vwire_39_17;
	reg signed[17:0] vreg_39_17;
	node n39_17(.left(vreg_38_17), .right(vreg_40_17), .up(vreg_39_18), .down(vreg_39_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_17), .sw(sw));
	wire signed[17:0] vwire_39_18;
	reg signed[17:0] vreg_39_18;
	node n39_18(.left(vreg_38_18), .right(vreg_40_18), .up(vreg_39_19), .down(vreg_39_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_18), .sw(sw));
	wire signed[17:0] vwire_39_19;
	reg signed[17:0] vreg_39_19;
	node n39_19(.left(vreg_38_19), .right(vreg_40_19), .up(vreg_39_20), .down(vreg_39_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_19), .sw(sw));
	wire signed[17:0] vwire_39_20;
	reg signed[17:0] vreg_39_20;
	node n39_20(.left(vreg_38_20), .right(vreg_40_20), .up(vreg_39_21), .down(vreg_39_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_20), .sw(sw));
	wire signed[17:0] vwire_39_21;
	reg signed[17:0] vreg_39_21;
	node n39_21(.left(vreg_38_21), .right(vreg_40_21), .up(vreg_39_22), .down(vreg_39_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_21), .sw(sw));
	wire signed[17:0] vwire_39_22;
	reg signed[17:0] vreg_39_22;
	node n39_22(.left(vreg_38_22), .right(vreg_40_22), .up(vreg_39_23), .down(vreg_39_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_22), .sw(sw));
	wire signed[17:0] vwire_39_23;
	reg signed[17:0] vreg_39_23;
	node n39_23(.left(vreg_38_23), .right(vreg_40_23), .up(vreg_39_24), .down(vreg_39_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_23), .sw(sw));
	wire signed[17:0] vwire_39_24;
	reg signed[17:0] vreg_39_24;
	node n39_24(.left(vreg_38_24), .right(vreg_40_24), .up(vreg_39_25), .down(vreg_39_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_24), .sw(sw));
	wire signed[17:0] vwire_39_25;
	reg signed[17:0] vreg_39_25;
	node n39_25(.left(vreg_38_25), .right(vreg_40_25), .up(vreg_39_26), .down(vreg_39_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_25), .sw(sw));
	wire signed[17:0] vwire_39_26;
	reg signed[17:0] vreg_39_26;
	node n39_26(.left(vreg_38_26), .right(vreg_40_26), .up(vreg_39_27), .down(vreg_39_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_26), .sw(sw));
	wire signed[17:0] vwire_39_27;
	reg signed[17:0] vreg_39_27;
	node n39_27(.left(vreg_38_27), .right(vreg_40_27), .up(vreg_39_28), .down(vreg_39_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_27), .sw(sw));
	wire signed[17:0] vwire_39_28;
	reg signed[17:0] vreg_39_28;
	node n39_28(.left(vreg_38_28), .right(vreg_40_28), .up(vreg_39_29), .down(vreg_39_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_28), .sw(sw));
	wire signed[17:0] vwire_39_29;
	reg signed[17:0] vreg_39_29;
	node n39_29(.left(vreg_38_29), .right(vreg_40_29), .up(vreg_39_30), .down(vreg_39_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_29), .sw(sw));
	wire signed[17:0] vwire_39_30;
	reg signed[17:0] vreg_39_30;
	node n39_30(.left(vreg_38_30), .right(vreg_40_30), .up(vreg_39_31), .down(vreg_39_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_30), .sw(sw));
	wire signed[17:0] vwire_39_31;
	reg signed[17:0] vreg_39_31;
	node n39_31(.left(vreg_38_31), .right(vreg_40_31), .up(vreg_39_32), .down(vreg_39_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_31), .sw(sw));
	wire signed[17:0] vwire_39_32;
	reg signed[17:0] vreg_39_32;
	node n39_32(.left(vreg_38_32), .right(vreg_40_32), .up(vreg_39_33), .down(vreg_39_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_32), .sw(sw));
	wire signed[17:0] vwire_39_33;
	reg signed[17:0] vreg_39_33;
	node n39_33(.left(vreg_38_33), .right(vreg_40_33), .up(vreg_39_34), .down(vreg_39_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_33), .sw(sw));
	wire signed[17:0] vwire_39_34;
	reg signed[17:0] vreg_39_34;
	node n39_34(.left(vreg_38_34), .right(vreg_40_34), .up(vreg_39_35), .down(vreg_39_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_34), .sw(sw));
	wire signed[17:0] vwire_39_35;
	reg signed[17:0] vreg_39_35;
	node n39_35(.left(vreg_38_35), .right(vreg_40_35), .up(vreg_39_36), .down(vreg_39_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_35), .sw(sw));
	wire signed[17:0] vwire_39_36;
	reg signed[17:0] vreg_39_36;
	node n39_36(.left(vreg_38_36), .right(vreg_40_36), .up(vreg_39_37), .down(vreg_39_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_36), .sw(sw));
	wire signed[17:0] vwire_39_37;
	reg signed[17:0] vreg_39_37;
	node n39_37(.left(vreg_38_37), .right(vreg_40_37), .up(vreg_39_38), .down(vreg_39_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_37), .sw(sw));
	wire signed[17:0] vwire_39_38;
	reg signed[17:0] vreg_39_38;
	node n39_38(.left(vreg_38_38), .right(vreg_40_38), .up(vreg_39_39), .down(vreg_39_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_38), .sw(sw));
	wire signed[17:0] vwire_39_39;
	reg signed[17:0] vreg_39_39;
	node n39_39(.left(vreg_38_39), .right(vreg_40_39), .up(vreg_39_40), .down(vreg_39_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_39), .sw(sw));
	wire signed[17:0] vwire_39_40;
	reg signed[17:0] vreg_39_40;
	node n39_40(.left(vreg_38_40), .right(vreg_40_40), .up(vreg_39_41), .down(vreg_39_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_40), .sw(sw));
	wire signed[17:0] vwire_39_41;
	reg signed[17:0] vreg_39_41;
	node n39_41(.left(vreg_38_41), .right(vreg_40_41), .up(vreg_39_42), .down(vreg_39_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_41), .sw(sw));
	wire signed[17:0] vwire_39_42;
	reg signed[17:0] vreg_39_42;
	node n39_42(.left(vreg_38_42), .right(vreg_40_42), .up(vreg_39_43), .down(vreg_39_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_42), .sw(sw));
	wire signed[17:0] vwire_39_43;
	reg signed[17:0] vreg_39_43;
	node n39_43(.left(vreg_38_43), .right(vreg_40_43), .up(vreg_39_44), .down(vreg_39_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_43), .sw(sw));
	wire signed[17:0] vwire_39_44;
	reg signed[17:0] vreg_39_44;
	node n39_44(.left(vreg_38_44), .right(vreg_40_44), .up(vreg_39_45), .down(vreg_39_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_44), .sw(sw));
	wire signed[17:0] vwire_39_45;
	reg signed[17:0] vreg_39_45;
	node n39_45(.left(vreg_38_45), .right(vreg_40_45), .up(vreg_39_46), .down(vreg_39_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_45), .sw(sw));
	wire signed[17:0] vwire_39_46;
	reg signed[17:0] vreg_39_46;
	node n39_46(.left(vreg_38_46), .right(vreg_40_46), .up(vreg_39_47), .down(vreg_39_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_46), .sw(sw));
	wire signed[17:0] vwire_39_47;
	reg signed[17:0] vreg_39_47;
	node n39_47(.left(vreg_38_47), .right(vreg_40_47), .up(vreg_39_48), .down(vreg_39_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_47), .sw(sw));
	wire signed[17:0] vwire_39_48;
	reg signed[17:0] vreg_39_48;
	node n39_48(.left(vreg_38_48), .right(vreg_40_48), .up(vreg_39_49), .down(vreg_39_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_48), .sw(sw));
	wire signed[17:0] vwire_39_49;
	reg signed[17:0] vreg_39_49;
	node n39_49(.left(vreg_38_49), .right(vreg_40_49), .up(18'b0), .down(vreg_39_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_39_49), .sw(sw));
	wire signed[17:0] vwire_40_0;
	reg signed[17:0] vreg_40_0;
	node n40_0(.left(vreg_39_0), .right(vreg_41_0), .up(vreg_40_1), .down(vreg_40_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_0), .sw(sw));
	wire signed[17:0] vwire_40_1;
	reg signed[17:0] vreg_40_1;
	node n40_1(.left(vreg_39_1), .right(vreg_41_1), .up(vreg_40_2), .down(vreg_40_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_1), .sw(sw));
	wire signed[17:0] vwire_40_2;
	reg signed[17:0] vreg_40_2;
	node n40_2(.left(vreg_39_2), .right(vreg_41_2), .up(vreg_40_3), .down(vreg_40_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_2), .sw(sw));
	wire signed[17:0] vwire_40_3;
	reg signed[17:0] vreg_40_3;
	node n40_3(.left(vreg_39_3), .right(vreg_41_3), .up(vreg_40_4), .down(vreg_40_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_3), .sw(sw));
	wire signed[17:0] vwire_40_4;
	reg signed[17:0] vreg_40_4;
	node n40_4(.left(vreg_39_4), .right(vreg_41_4), .up(vreg_40_5), .down(vreg_40_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_4), .sw(sw));
	wire signed[17:0] vwire_40_5;
	reg signed[17:0] vreg_40_5;
	node n40_5(.left(vreg_39_5), .right(vreg_41_5), .up(vreg_40_6), .down(vreg_40_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_5), .sw(sw));
	wire signed[17:0] vwire_40_6;
	reg signed[17:0] vreg_40_6;
	node n40_6(.left(vreg_39_6), .right(vreg_41_6), .up(vreg_40_7), .down(vreg_40_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_6), .sw(sw));
	wire signed[17:0] vwire_40_7;
	reg signed[17:0] vreg_40_7;
	node n40_7(.left(vreg_39_7), .right(vreg_41_7), .up(vreg_40_8), .down(vreg_40_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_7), .sw(sw));
	wire signed[17:0] vwire_40_8;
	reg signed[17:0] vreg_40_8;
	node n40_8(.left(vreg_39_8), .right(vreg_41_8), .up(vreg_40_9), .down(vreg_40_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_8), .sw(sw));
	wire signed[17:0] vwire_40_9;
	reg signed[17:0] vreg_40_9;
	node n40_9(.left(vreg_39_9), .right(vreg_41_9), .up(vreg_40_10), .down(vreg_40_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_9), .sw(sw));
	wire signed[17:0] vwire_40_10;
	reg signed[17:0] vreg_40_10;
	node n40_10(.left(vreg_39_10), .right(vreg_41_10), .up(vreg_40_11), .down(vreg_40_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_10), .sw(sw));
	wire signed[17:0] vwire_40_11;
	reg signed[17:0] vreg_40_11;
	node n40_11(.left(vreg_39_11), .right(vreg_41_11), .up(vreg_40_12), .down(vreg_40_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_11), .sw(sw));
	wire signed[17:0] vwire_40_12;
	reg signed[17:0] vreg_40_12;
	node n40_12(.left(vreg_39_12), .right(vreg_41_12), .up(vreg_40_13), .down(vreg_40_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_12), .sw(sw));
	wire signed[17:0] vwire_40_13;
	reg signed[17:0] vreg_40_13;
	node n40_13(.left(vreg_39_13), .right(vreg_41_13), .up(vreg_40_14), .down(vreg_40_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_13), .sw(sw));
	wire signed[17:0] vwire_40_14;
	reg signed[17:0] vreg_40_14;
	node n40_14(.left(vreg_39_14), .right(vreg_41_14), .up(vreg_40_15), .down(vreg_40_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_14), .sw(sw));
	wire signed[17:0] vwire_40_15;
	reg signed[17:0] vreg_40_15;
	node n40_15(.left(vreg_39_15), .right(vreg_41_15), .up(vreg_40_16), .down(vreg_40_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_15), .sw(sw));
	wire signed[17:0] vwire_40_16;
	reg signed[17:0] vreg_40_16;
	node n40_16(.left(vreg_39_16), .right(vreg_41_16), .up(vreg_40_17), .down(vreg_40_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_16), .sw(sw));
	wire signed[17:0] vwire_40_17;
	reg signed[17:0] vreg_40_17;
	node n40_17(.left(vreg_39_17), .right(vreg_41_17), .up(vreg_40_18), .down(vreg_40_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_17), .sw(sw));
	wire signed[17:0] vwire_40_18;
	reg signed[17:0] vreg_40_18;
	node n40_18(.left(vreg_39_18), .right(vreg_41_18), .up(vreg_40_19), .down(vreg_40_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_18), .sw(sw));
	wire signed[17:0] vwire_40_19;
	reg signed[17:0] vreg_40_19;
	node n40_19(.left(vreg_39_19), .right(vreg_41_19), .up(vreg_40_20), .down(vreg_40_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_19), .sw(sw));
	wire signed[17:0] vwire_40_20;
	reg signed[17:0] vreg_40_20;
	node n40_20(.left(vreg_39_20), .right(vreg_41_20), .up(vreg_40_21), .down(vreg_40_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_20), .sw(sw));
	wire signed[17:0] vwire_40_21;
	reg signed[17:0] vreg_40_21;
	node n40_21(.left(vreg_39_21), .right(vreg_41_21), .up(vreg_40_22), .down(vreg_40_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_21), .sw(sw));
	wire signed[17:0] vwire_40_22;
	reg signed[17:0] vreg_40_22;
	node n40_22(.left(vreg_39_22), .right(vreg_41_22), .up(vreg_40_23), .down(vreg_40_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_22), .sw(sw));
	wire signed[17:0] vwire_40_23;
	reg signed[17:0] vreg_40_23;
	node n40_23(.left(vreg_39_23), .right(vreg_41_23), .up(vreg_40_24), .down(vreg_40_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_23), .sw(sw));
	wire signed[17:0] vwire_40_24;
	reg signed[17:0] vreg_40_24;
	node n40_24(.left(vreg_39_24), .right(vreg_41_24), .up(vreg_40_25), .down(vreg_40_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_24), .sw(sw));
	wire signed[17:0] vwire_40_25;
	reg signed[17:0] vreg_40_25;
	node n40_25(.left(vreg_39_25), .right(vreg_41_25), .up(vreg_40_26), .down(vreg_40_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_25), .sw(sw));
	wire signed[17:0] vwire_40_26;
	reg signed[17:0] vreg_40_26;
	node n40_26(.left(vreg_39_26), .right(vreg_41_26), .up(vreg_40_27), .down(vreg_40_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_26), .sw(sw));
	wire signed[17:0] vwire_40_27;
	reg signed[17:0] vreg_40_27;
	node n40_27(.left(vreg_39_27), .right(vreg_41_27), .up(vreg_40_28), .down(vreg_40_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_27), .sw(sw));
	wire signed[17:0] vwire_40_28;
	reg signed[17:0] vreg_40_28;
	node n40_28(.left(vreg_39_28), .right(vreg_41_28), .up(vreg_40_29), .down(vreg_40_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_28), .sw(sw));
	wire signed[17:0] vwire_40_29;
	reg signed[17:0] vreg_40_29;
	node n40_29(.left(vreg_39_29), .right(vreg_41_29), .up(vreg_40_30), .down(vreg_40_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_29), .sw(sw));
	wire signed[17:0] vwire_40_30;
	reg signed[17:0] vreg_40_30;
	node n40_30(.left(vreg_39_30), .right(vreg_41_30), .up(vreg_40_31), .down(vreg_40_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_30), .sw(sw));
	wire signed[17:0] vwire_40_31;
	reg signed[17:0] vreg_40_31;
	node n40_31(.left(vreg_39_31), .right(vreg_41_31), .up(vreg_40_32), .down(vreg_40_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_31), .sw(sw));
	wire signed[17:0] vwire_40_32;
	reg signed[17:0] vreg_40_32;
	node n40_32(.left(vreg_39_32), .right(vreg_41_32), .up(vreg_40_33), .down(vreg_40_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_32), .sw(sw));
	wire signed[17:0] vwire_40_33;
	reg signed[17:0] vreg_40_33;
	node n40_33(.left(vreg_39_33), .right(vreg_41_33), .up(vreg_40_34), .down(vreg_40_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_33), .sw(sw));
	wire signed[17:0] vwire_40_34;
	reg signed[17:0] vreg_40_34;
	node n40_34(.left(vreg_39_34), .right(vreg_41_34), .up(vreg_40_35), .down(vreg_40_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_34), .sw(sw));
	wire signed[17:0] vwire_40_35;
	reg signed[17:0] vreg_40_35;
	node n40_35(.left(vreg_39_35), .right(vreg_41_35), .up(vreg_40_36), .down(vreg_40_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_35), .sw(sw));
	wire signed[17:0] vwire_40_36;
	reg signed[17:0] vreg_40_36;
	node n40_36(.left(vreg_39_36), .right(vreg_41_36), .up(vreg_40_37), .down(vreg_40_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_36), .sw(sw));
	wire signed[17:0] vwire_40_37;
	reg signed[17:0] vreg_40_37;
	node n40_37(.left(vreg_39_37), .right(vreg_41_37), .up(vreg_40_38), .down(vreg_40_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_37), .sw(sw));
	wire signed[17:0] vwire_40_38;
	reg signed[17:0] vreg_40_38;
	node n40_38(.left(vreg_39_38), .right(vreg_41_38), .up(vreg_40_39), .down(vreg_40_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_38), .sw(sw));
	wire signed[17:0] vwire_40_39;
	reg signed[17:0] vreg_40_39;
	node n40_39(.left(vreg_39_39), .right(vreg_41_39), .up(vreg_40_40), .down(vreg_40_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_39), .sw(sw));
	wire signed[17:0] vwire_40_40;
	reg signed[17:0] vreg_40_40;
	node n40_40(.left(vreg_39_40), .right(vreg_41_40), .up(vreg_40_41), .down(vreg_40_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_40), .sw(sw));
	wire signed[17:0] vwire_40_41;
	reg signed[17:0] vreg_40_41;
	node n40_41(.left(vreg_39_41), .right(vreg_41_41), .up(vreg_40_42), .down(vreg_40_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_41), .sw(sw));
	wire signed[17:0] vwire_40_42;
	reg signed[17:0] vreg_40_42;
	node n40_42(.left(vreg_39_42), .right(vreg_41_42), .up(vreg_40_43), .down(vreg_40_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_42), .sw(sw));
	wire signed[17:0] vwire_40_43;
	reg signed[17:0] vreg_40_43;
	node n40_43(.left(vreg_39_43), .right(vreg_41_43), .up(vreg_40_44), .down(vreg_40_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_43), .sw(sw));
	wire signed[17:0] vwire_40_44;
	reg signed[17:0] vreg_40_44;
	node n40_44(.left(vreg_39_44), .right(vreg_41_44), .up(vreg_40_45), .down(vreg_40_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_44), .sw(sw));
	wire signed[17:0] vwire_40_45;
	reg signed[17:0] vreg_40_45;
	node n40_45(.left(vreg_39_45), .right(vreg_41_45), .up(vreg_40_46), .down(vreg_40_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_45), .sw(sw));
	wire signed[17:0] vwire_40_46;
	reg signed[17:0] vreg_40_46;
	node n40_46(.left(vreg_39_46), .right(vreg_41_46), .up(vreg_40_47), .down(vreg_40_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_46), .sw(sw));
	wire signed[17:0] vwire_40_47;
	reg signed[17:0] vreg_40_47;
	node n40_47(.left(vreg_39_47), .right(vreg_41_47), .up(vreg_40_48), .down(vreg_40_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_47), .sw(sw));
	wire signed[17:0] vwire_40_48;
	reg signed[17:0] vreg_40_48;
	node n40_48(.left(vreg_39_48), .right(vreg_41_48), .up(vreg_40_49), .down(vreg_40_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_48), .sw(sw));
	wire signed[17:0] vwire_40_49;
	reg signed[17:0] vreg_40_49;
	node n40_49(.left(vreg_39_49), .right(vreg_41_49), .up(18'b0), .down(vreg_40_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_40_49), .sw(sw));
	wire signed[17:0] vwire_41_0;
	reg signed[17:0] vreg_41_0;
	node n41_0(.left(vreg_40_0), .right(vreg_42_0), .up(vreg_41_1), .down(vreg_41_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_0), .sw(sw));
	wire signed[17:0] vwire_41_1;
	reg signed[17:0] vreg_41_1;
	node n41_1(.left(vreg_40_1), .right(vreg_42_1), .up(vreg_41_2), .down(vreg_41_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_1), .sw(sw));
	wire signed[17:0] vwire_41_2;
	reg signed[17:0] vreg_41_2;
	node n41_2(.left(vreg_40_2), .right(vreg_42_2), .up(vreg_41_3), .down(vreg_41_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_2), .sw(sw));
	wire signed[17:0] vwire_41_3;
	reg signed[17:0] vreg_41_3;
	node n41_3(.left(vreg_40_3), .right(vreg_42_3), .up(vreg_41_4), .down(vreg_41_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_3), .sw(sw));
	wire signed[17:0] vwire_41_4;
	reg signed[17:0] vreg_41_4;
	node n41_4(.left(vreg_40_4), .right(vreg_42_4), .up(vreg_41_5), .down(vreg_41_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_4), .sw(sw));
	wire signed[17:0] vwire_41_5;
	reg signed[17:0] vreg_41_5;
	node n41_5(.left(vreg_40_5), .right(vreg_42_5), .up(vreg_41_6), .down(vreg_41_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_5), .sw(sw));
	wire signed[17:0] vwire_41_6;
	reg signed[17:0] vreg_41_6;
	node n41_6(.left(vreg_40_6), .right(vreg_42_6), .up(vreg_41_7), .down(vreg_41_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_6), .sw(sw));
	wire signed[17:0] vwire_41_7;
	reg signed[17:0] vreg_41_7;
	node n41_7(.left(vreg_40_7), .right(vreg_42_7), .up(vreg_41_8), .down(vreg_41_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_7), .sw(sw));
	wire signed[17:0] vwire_41_8;
	reg signed[17:0] vreg_41_8;
	node n41_8(.left(vreg_40_8), .right(vreg_42_8), .up(vreg_41_9), .down(vreg_41_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_8), .sw(sw));
	wire signed[17:0] vwire_41_9;
	reg signed[17:0] vreg_41_9;
	node n41_9(.left(vreg_40_9), .right(vreg_42_9), .up(vreg_41_10), .down(vreg_41_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_9), .sw(sw));
	wire signed[17:0] vwire_41_10;
	reg signed[17:0] vreg_41_10;
	node n41_10(.left(vreg_40_10), .right(vreg_42_10), .up(vreg_41_11), .down(vreg_41_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_10), .sw(sw));
	wire signed[17:0] vwire_41_11;
	reg signed[17:0] vreg_41_11;
	node n41_11(.left(vreg_40_11), .right(vreg_42_11), .up(vreg_41_12), .down(vreg_41_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_11), .sw(sw));
	wire signed[17:0] vwire_41_12;
	reg signed[17:0] vreg_41_12;
	node n41_12(.left(vreg_40_12), .right(vreg_42_12), .up(vreg_41_13), .down(vreg_41_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_12), .sw(sw));
	wire signed[17:0] vwire_41_13;
	reg signed[17:0] vreg_41_13;
	node n41_13(.left(vreg_40_13), .right(vreg_42_13), .up(vreg_41_14), .down(vreg_41_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_13), .sw(sw));
	wire signed[17:0] vwire_41_14;
	reg signed[17:0] vreg_41_14;
	node n41_14(.left(vreg_40_14), .right(vreg_42_14), .up(vreg_41_15), .down(vreg_41_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_14), .sw(sw));
	wire signed[17:0] vwire_41_15;
	reg signed[17:0] vreg_41_15;
	node n41_15(.left(vreg_40_15), .right(vreg_42_15), .up(vreg_41_16), .down(vreg_41_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_15), .sw(sw));
	wire signed[17:0] vwire_41_16;
	reg signed[17:0] vreg_41_16;
	node n41_16(.left(vreg_40_16), .right(vreg_42_16), .up(vreg_41_17), .down(vreg_41_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_16), .sw(sw));
	wire signed[17:0] vwire_41_17;
	reg signed[17:0] vreg_41_17;
	node n41_17(.left(vreg_40_17), .right(vreg_42_17), .up(vreg_41_18), .down(vreg_41_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_17), .sw(sw));
	wire signed[17:0] vwire_41_18;
	reg signed[17:0] vreg_41_18;
	node n41_18(.left(vreg_40_18), .right(vreg_42_18), .up(vreg_41_19), .down(vreg_41_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_18), .sw(sw));
	wire signed[17:0] vwire_41_19;
	reg signed[17:0] vreg_41_19;
	node n41_19(.left(vreg_40_19), .right(vreg_42_19), .up(vreg_41_20), .down(vreg_41_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_19), .sw(sw));
	wire signed[17:0] vwire_41_20;
	reg signed[17:0] vreg_41_20;
	node n41_20(.left(vreg_40_20), .right(vreg_42_20), .up(vreg_41_21), .down(vreg_41_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_20), .sw(sw));
	wire signed[17:0] vwire_41_21;
	reg signed[17:0] vreg_41_21;
	node n41_21(.left(vreg_40_21), .right(vreg_42_21), .up(vreg_41_22), .down(vreg_41_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_21), .sw(sw));
	wire signed[17:0] vwire_41_22;
	reg signed[17:0] vreg_41_22;
	node n41_22(.left(vreg_40_22), .right(vreg_42_22), .up(vreg_41_23), .down(vreg_41_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_22), .sw(sw));
	wire signed[17:0] vwire_41_23;
	reg signed[17:0] vreg_41_23;
	node n41_23(.left(vreg_40_23), .right(vreg_42_23), .up(vreg_41_24), .down(vreg_41_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_23), .sw(sw));
	wire signed[17:0] vwire_41_24;
	reg signed[17:0] vreg_41_24;
	node n41_24(.left(vreg_40_24), .right(vreg_42_24), .up(vreg_41_25), .down(vreg_41_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_24), .sw(sw));
	wire signed[17:0] vwire_41_25;
	reg signed[17:0] vreg_41_25;
	node n41_25(.left(vreg_40_25), .right(vreg_42_25), .up(vreg_41_26), .down(vreg_41_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_25), .sw(sw));
	wire signed[17:0] vwire_41_26;
	reg signed[17:0] vreg_41_26;
	node n41_26(.left(vreg_40_26), .right(vreg_42_26), .up(vreg_41_27), .down(vreg_41_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_26), .sw(sw));
	wire signed[17:0] vwire_41_27;
	reg signed[17:0] vreg_41_27;
	node n41_27(.left(vreg_40_27), .right(vreg_42_27), .up(vreg_41_28), .down(vreg_41_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_27), .sw(sw));
	wire signed[17:0] vwire_41_28;
	reg signed[17:0] vreg_41_28;
	node n41_28(.left(vreg_40_28), .right(vreg_42_28), .up(vreg_41_29), .down(vreg_41_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_28), .sw(sw));
	wire signed[17:0] vwire_41_29;
	reg signed[17:0] vreg_41_29;
	node n41_29(.left(vreg_40_29), .right(vreg_42_29), .up(vreg_41_30), .down(vreg_41_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_29), .sw(sw));
	wire signed[17:0] vwire_41_30;
	reg signed[17:0] vreg_41_30;
	node n41_30(.left(vreg_40_30), .right(vreg_42_30), .up(vreg_41_31), .down(vreg_41_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_30), .sw(sw));
	wire signed[17:0] vwire_41_31;
	reg signed[17:0] vreg_41_31;
	node n41_31(.left(vreg_40_31), .right(vreg_42_31), .up(vreg_41_32), .down(vreg_41_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_31), .sw(sw));
	wire signed[17:0] vwire_41_32;
	reg signed[17:0] vreg_41_32;
	node n41_32(.left(vreg_40_32), .right(vreg_42_32), .up(vreg_41_33), .down(vreg_41_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_32), .sw(sw));
	wire signed[17:0] vwire_41_33;
	reg signed[17:0] vreg_41_33;
	node n41_33(.left(vreg_40_33), .right(vreg_42_33), .up(vreg_41_34), .down(vreg_41_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_33), .sw(sw));
	wire signed[17:0] vwire_41_34;
	reg signed[17:0] vreg_41_34;
	node n41_34(.left(vreg_40_34), .right(vreg_42_34), .up(vreg_41_35), .down(vreg_41_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_34), .sw(sw));
	wire signed[17:0] vwire_41_35;
	reg signed[17:0] vreg_41_35;
	node n41_35(.left(vreg_40_35), .right(vreg_42_35), .up(vreg_41_36), .down(vreg_41_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_35), .sw(sw));
	wire signed[17:0] vwire_41_36;
	reg signed[17:0] vreg_41_36;
	node n41_36(.left(vreg_40_36), .right(vreg_42_36), .up(vreg_41_37), .down(vreg_41_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_36), .sw(sw));
	wire signed[17:0] vwire_41_37;
	reg signed[17:0] vreg_41_37;
	node n41_37(.left(vreg_40_37), .right(vreg_42_37), .up(vreg_41_38), .down(vreg_41_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_37), .sw(sw));
	wire signed[17:0] vwire_41_38;
	reg signed[17:0] vreg_41_38;
	node n41_38(.left(vreg_40_38), .right(vreg_42_38), .up(vreg_41_39), .down(vreg_41_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_38), .sw(sw));
	wire signed[17:0] vwire_41_39;
	reg signed[17:0] vreg_41_39;
	node n41_39(.left(vreg_40_39), .right(vreg_42_39), .up(vreg_41_40), .down(vreg_41_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_39), .sw(sw));
	wire signed[17:0] vwire_41_40;
	reg signed[17:0] vreg_41_40;
	node n41_40(.left(vreg_40_40), .right(vreg_42_40), .up(vreg_41_41), .down(vreg_41_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_40), .sw(sw));
	wire signed[17:0] vwire_41_41;
	reg signed[17:0] vreg_41_41;
	node n41_41(.left(vreg_40_41), .right(vreg_42_41), .up(vreg_41_42), .down(vreg_41_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_41), .sw(sw));
	wire signed[17:0] vwire_41_42;
	reg signed[17:0] vreg_41_42;
	node n41_42(.left(vreg_40_42), .right(vreg_42_42), .up(vreg_41_43), .down(vreg_41_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_42), .sw(sw));
	wire signed[17:0] vwire_41_43;
	reg signed[17:0] vreg_41_43;
	node n41_43(.left(vreg_40_43), .right(vreg_42_43), .up(vreg_41_44), .down(vreg_41_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_43), .sw(sw));
	wire signed[17:0] vwire_41_44;
	reg signed[17:0] vreg_41_44;
	node n41_44(.left(vreg_40_44), .right(vreg_42_44), .up(vreg_41_45), .down(vreg_41_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_44), .sw(sw));
	wire signed[17:0] vwire_41_45;
	reg signed[17:0] vreg_41_45;
	node n41_45(.left(vreg_40_45), .right(vreg_42_45), .up(vreg_41_46), .down(vreg_41_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_45), .sw(sw));
	wire signed[17:0] vwire_41_46;
	reg signed[17:0] vreg_41_46;
	node n41_46(.left(vreg_40_46), .right(vreg_42_46), .up(vreg_41_47), .down(vreg_41_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_46), .sw(sw));
	wire signed[17:0] vwire_41_47;
	reg signed[17:0] vreg_41_47;
	node n41_47(.left(vreg_40_47), .right(vreg_42_47), .up(vreg_41_48), .down(vreg_41_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_47), .sw(sw));
	wire signed[17:0] vwire_41_48;
	reg signed[17:0] vreg_41_48;
	node n41_48(.left(vreg_40_48), .right(vreg_42_48), .up(vreg_41_49), .down(vreg_41_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_48), .sw(sw));
	wire signed[17:0] vwire_41_49;
	reg signed[17:0] vreg_41_49;
	node n41_49(.left(vreg_40_49), .right(vreg_42_49), .up(18'b0), .down(vreg_41_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_41_49), .sw(sw));
	wire signed[17:0] vwire_42_0;
	reg signed[17:0] vreg_42_0;
	node n42_0(.left(vreg_41_0), .right(vreg_43_0), .up(vreg_42_1), .down(vreg_42_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_0), .sw(sw));
	wire signed[17:0] vwire_42_1;
	reg signed[17:0] vreg_42_1;
	node n42_1(.left(vreg_41_1), .right(vreg_43_1), .up(vreg_42_2), .down(vreg_42_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_1), .sw(sw));
	wire signed[17:0] vwire_42_2;
	reg signed[17:0] vreg_42_2;
	node n42_2(.left(vreg_41_2), .right(vreg_43_2), .up(vreg_42_3), .down(vreg_42_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_2), .sw(sw));
	wire signed[17:0] vwire_42_3;
	reg signed[17:0] vreg_42_3;
	node n42_3(.left(vreg_41_3), .right(vreg_43_3), .up(vreg_42_4), .down(vreg_42_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_3), .sw(sw));
	wire signed[17:0] vwire_42_4;
	reg signed[17:0] vreg_42_4;
	node n42_4(.left(vreg_41_4), .right(vreg_43_4), .up(vreg_42_5), .down(vreg_42_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_4), .sw(sw));
	wire signed[17:0] vwire_42_5;
	reg signed[17:0] vreg_42_5;
	node n42_5(.left(vreg_41_5), .right(vreg_43_5), .up(vreg_42_6), .down(vreg_42_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_5), .sw(sw));
	wire signed[17:0] vwire_42_6;
	reg signed[17:0] vreg_42_6;
	node n42_6(.left(vreg_41_6), .right(vreg_43_6), .up(vreg_42_7), .down(vreg_42_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_6), .sw(sw));
	wire signed[17:0] vwire_42_7;
	reg signed[17:0] vreg_42_7;
	node n42_7(.left(vreg_41_7), .right(vreg_43_7), .up(vreg_42_8), .down(vreg_42_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_7), .sw(sw));
	wire signed[17:0] vwire_42_8;
	reg signed[17:0] vreg_42_8;
	node n42_8(.left(vreg_41_8), .right(vreg_43_8), .up(vreg_42_9), .down(vreg_42_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_8), .sw(sw));
	wire signed[17:0] vwire_42_9;
	reg signed[17:0] vreg_42_9;
	node n42_9(.left(vreg_41_9), .right(vreg_43_9), .up(vreg_42_10), .down(vreg_42_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_9), .sw(sw));
	wire signed[17:0] vwire_42_10;
	reg signed[17:0] vreg_42_10;
	node n42_10(.left(vreg_41_10), .right(vreg_43_10), .up(vreg_42_11), .down(vreg_42_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_10), .sw(sw));
	wire signed[17:0] vwire_42_11;
	reg signed[17:0] vreg_42_11;
	node n42_11(.left(vreg_41_11), .right(vreg_43_11), .up(vreg_42_12), .down(vreg_42_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_11), .sw(sw));
	wire signed[17:0] vwire_42_12;
	reg signed[17:0] vreg_42_12;
	node n42_12(.left(vreg_41_12), .right(vreg_43_12), .up(vreg_42_13), .down(vreg_42_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_12), .sw(sw));
	wire signed[17:0] vwire_42_13;
	reg signed[17:0] vreg_42_13;
	node n42_13(.left(vreg_41_13), .right(vreg_43_13), .up(vreg_42_14), .down(vreg_42_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_13), .sw(sw));
	wire signed[17:0] vwire_42_14;
	reg signed[17:0] vreg_42_14;
	node n42_14(.left(vreg_41_14), .right(vreg_43_14), .up(vreg_42_15), .down(vreg_42_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_14), .sw(sw));
	wire signed[17:0] vwire_42_15;
	reg signed[17:0] vreg_42_15;
	node n42_15(.left(vreg_41_15), .right(vreg_43_15), .up(vreg_42_16), .down(vreg_42_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_15), .sw(sw));
	wire signed[17:0] vwire_42_16;
	reg signed[17:0] vreg_42_16;
	node n42_16(.left(vreg_41_16), .right(vreg_43_16), .up(vreg_42_17), .down(vreg_42_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_16), .sw(sw));
	wire signed[17:0] vwire_42_17;
	reg signed[17:0] vreg_42_17;
	node n42_17(.left(vreg_41_17), .right(vreg_43_17), .up(vreg_42_18), .down(vreg_42_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_17), .sw(sw));
	wire signed[17:0] vwire_42_18;
	reg signed[17:0] vreg_42_18;
	node n42_18(.left(vreg_41_18), .right(vreg_43_18), .up(vreg_42_19), .down(vreg_42_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_18), .sw(sw));
	wire signed[17:0] vwire_42_19;
	reg signed[17:0] vreg_42_19;
	node n42_19(.left(vreg_41_19), .right(vreg_43_19), .up(vreg_42_20), .down(vreg_42_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_19), .sw(sw));
	wire signed[17:0] vwire_42_20;
	reg signed[17:0] vreg_42_20;
	node n42_20(.left(vreg_41_20), .right(vreg_43_20), .up(vreg_42_21), .down(vreg_42_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_20), .sw(sw));
	wire signed[17:0] vwire_42_21;
	reg signed[17:0] vreg_42_21;
	node n42_21(.left(vreg_41_21), .right(vreg_43_21), .up(vreg_42_22), .down(vreg_42_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_21), .sw(sw));
	wire signed[17:0] vwire_42_22;
	reg signed[17:0] vreg_42_22;
	node n42_22(.left(vreg_41_22), .right(vreg_43_22), .up(vreg_42_23), .down(vreg_42_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_22), .sw(sw));
	wire signed[17:0] vwire_42_23;
	reg signed[17:0] vreg_42_23;
	node n42_23(.left(vreg_41_23), .right(vreg_43_23), .up(vreg_42_24), .down(vreg_42_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_23), .sw(sw));
	wire signed[17:0] vwire_42_24;
	reg signed[17:0] vreg_42_24;
	node n42_24(.left(vreg_41_24), .right(vreg_43_24), .up(vreg_42_25), .down(vreg_42_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_24), .sw(sw));
	wire signed[17:0] vwire_42_25;
	reg signed[17:0] vreg_42_25;
	node n42_25(.left(vreg_41_25), .right(vreg_43_25), .up(vreg_42_26), .down(vreg_42_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_25), .sw(sw));
	wire signed[17:0] vwire_42_26;
	reg signed[17:0] vreg_42_26;
	node n42_26(.left(vreg_41_26), .right(vreg_43_26), .up(vreg_42_27), .down(vreg_42_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_26), .sw(sw));
	wire signed[17:0] vwire_42_27;
	reg signed[17:0] vreg_42_27;
	node n42_27(.left(vreg_41_27), .right(vreg_43_27), .up(vreg_42_28), .down(vreg_42_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_27), .sw(sw));
	wire signed[17:0] vwire_42_28;
	reg signed[17:0] vreg_42_28;
	node n42_28(.left(vreg_41_28), .right(vreg_43_28), .up(vreg_42_29), .down(vreg_42_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_28), .sw(sw));
	wire signed[17:0] vwire_42_29;
	reg signed[17:0] vreg_42_29;
	node n42_29(.left(vreg_41_29), .right(vreg_43_29), .up(vreg_42_30), .down(vreg_42_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_29), .sw(sw));
	wire signed[17:0] vwire_42_30;
	reg signed[17:0] vreg_42_30;
	node n42_30(.left(vreg_41_30), .right(vreg_43_30), .up(vreg_42_31), .down(vreg_42_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_30), .sw(sw));
	wire signed[17:0] vwire_42_31;
	reg signed[17:0] vreg_42_31;
	node n42_31(.left(vreg_41_31), .right(vreg_43_31), .up(vreg_42_32), .down(vreg_42_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_31), .sw(sw));
	wire signed[17:0] vwire_42_32;
	reg signed[17:0] vreg_42_32;
	node n42_32(.left(vreg_41_32), .right(vreg_43_32), .up(vreg_42_33), .down(vreg_42_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_32), .sw(sw));
	wire signed[17:0] vwire_42_33;
	reg signed[17:0] vreg_42_33;
	node n42_33(.left(vreg_41_33), .right(vreg_43_33), .up(vreg_42_34), .down(vreg_42_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_33), .sw(sw));
	wire signed[17:0] vwire_42_34;
	reg signed[17:0] vreg_42_34;
	node n42_34(.left(vreg_41_34), .right(vreg_43_34), .up(vreg_42_35), .down(vreg_42_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_34), .sw(sw));
	wire signed[17:0] vwire_42_35;
	reg signed[17:0] vreg_42_35;
	node n42_35(.left(vreg_41_35), .right(vreg_43_35), .up(vreg_42_36), .down(vreg_42_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_35), .sw(sw));
	wire signed[17:0] vwire_42_36;
	reg signed[17:0] vreg_42_36;
	node n42_36(.left(vreg_41_36), .right(vreg_43_36), .up(vreg_42_37), .down(vreg_42_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_36), .sw(sw));
	wire signed[17:0] vwire_42_37;
	reg signed[17:0] vreg_42_37;
	node n42_37(.left(vreg_41_37), .right(vreg_43_37), .up(vreg_42_38), .down(vreg_42_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_37), .sw(sw));
	wire signed[17:0] vwire_42_38;
	reg signed[17:0] vreg_42_38;
	node n42_38(.left(vreg_41_38), .right(vreg_43_38), .up(vreg_42_39), .down(vreg_42_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_38), .sw(sw));
	wire signed[17:0] vwire_42_39;
	reg signed[17:0] vreg_42_39;
	node n42_39(.left(vreg_41_39), .right(vreg_43_39), .up(vreg_42_40), .down(vreg_42_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_39), .sw(sw));
	wire signed[17:0] vwire_42_40;
	reg signed[17:0] vreg_42_40;
	node n42_40(.left(vreg_41_40), .right(vreg_43_40), .up(vreg_42_41), .down(vreg_42_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_40), .sw(sw));
	wire signed[17:0] vwire_42_41;
	reg signed[17:0] vreg_42_41;
	node n42_41(.left(vreg_41_41), .right(vreg_43_41), .up(vreg_42_42), .down(vreg_42_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_41), .sw(sw));
	wire signed[17:0] vwire_42_42;
	reg signed[17:0] vreg_42_42;
	node n42_42(.left(vreg_41_42), .right(vreg_43_42), .up(vreg_42_43), .down(vreg_42_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_42), .sw(sw));
	wire signed[17:0] vwire_42_43;
	reg signed[17:0] vreg_42_43;
	node n42_43(.left(vreg_41_43), .right(vreg_43_43), .up(vreg_42_44), .down(vreg_42_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_43), .sw(sw));
	wire signed[17:0] vwire_42_44;
	reg signed[17:0] vreg_42_44;
	node n42_44(.left(vreg_41_44), .right(vreg_43_44), .up(vreg_42_45), .down(vreg_42_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_44), .sw(sw));
	wire signed[17:0] vwire_42_45;
	reg signed[17:0] vreg_42_45;
	node n42_45(.left(vreg_41_45), .right(vreg_43_45), .up(vreg_42_46), .down(vreg_42_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_45), .sw(sw));
	wire signed[17:0] vwire_42_46;
	reg signed[17:0] vreg_42_46;
	node n42_46(.left(vreg_41_46), .right(vreg_43_46), .up(vreg_42_47), .down(vreg_42_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_46), .sw(sw));
	wire signed[17:0] vwire_42_47;
	reg signed[17:0] vreg_42_47;
	node n42_47(.left(vreg_41_47), .right(vreg_43_47), .up(vreg_42_48), .down(vreg_42_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_47), .sw(sw));
	wire signed[17:0] vwire_42_48;
	reg signed[17:0] vreg_42_48;
	node n42_48(.left(vreg_41_48), .right(vreg_43_48), .up(vreg_42_49), .down(vreg_42_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_48), .sw(sw));
	wire signed[17:0] vwire_42_49;
	reg signed[17:0] vreg_42_49;
	node n42_49(.left(vreg_41_49), .right(vreg_43_49), .up(18'b0), .down(vreg_42_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_42_49), .sw(sw));
	wire signed[17:0] vwire_43_0;
	reg signed[17:0] vreg_43_0;
	node n43_0(.left(vreg_42_0), .right(vreg_44_0), .up(vreg_43_1), .down(vreg_43_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_0), .sw(sw));
	wire signed[17:0] vwire_43_1;
	reg signed[17:0] vreg_43_1;
	node n43_1(.left(vreg_42_1), .right(vreg_44_1), .up(vreg_43_2), .down(vreg_43_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_1), .sw(sw));
	wire signed[17:0] vwire_43_2;
	reg signed[17:0] vreg_43_2;
	node n43_2(.left(vreg_42_2), .right(vreg_44_2), .up(vreg_43_3), .down(vreg_43_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_2), .sw(sw));
	wire signed[17:0] vwire_43_3;
	reg signed[17:0] vreg_43_3;
	node n43_3(.left(vreg_42_3), .right(vreg_44_3), .up(vreg_43_4), .down(vreg_43_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_3), .sw(sw));
	wire signed[17:0] vwire_43_4;
	reg signed[17:0] vreg_43_4;
	node n43_4(.left(vreg_42_4), .right(vreg_44_4), .up(vreg_43_5), .down(vreg_43_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_4), .sw(sw));
	wire signed[17:0] vwire_43_5;
	reg signed[17:0] vreg_43_5;
	node n43_5(.left(vreg_42_5), .right(vreg_44_5), .up(vreg_43_6), .down(vreg_43_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_5), .sw(sw));
	wire signed[17:0] vwire_43_6;
	reg signed[17:0] vreg_43_6;
	node n43_6(.left(vreg_42_6), .right(vreg_44_6), .up(vreg_43_7), .down(vreg_43_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_6), .sw(sw));
	wire signed[17:0] vwire_43_7;
	reg signed[17:0] vreg_43_7;
	node n43_7(.left(vreg_42_7), .right(vreg_44_7), .up(vreg_43_8), .down(vreg_43_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_7), .sw(sw));
	wire signed[17:0] vwire_43_8;
	reg signed[17:0] vreg_43_8;
	node n43_8(.left(vreg_42_8), .right(vreg_44_8), .up(vreg_43_9), .down(vreg_43_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_8), .sw(sw));
	wire signed[17:0] vwire_43_9;
	reg signed[17:0] vreg_43_9;
	node n43_9(.left(vreg_42_9), .right(vreg_44_9), .up(vreg_43_10), .down(vreg_43_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_9), .sw(sw));
	wire signed[17:0] vwire_43_10;
	reg signed[17:0] vreg_43_10;
	node n43_10(.left(vreg_42_10), .right(vreg_44_10), .up(vreg_43_11), .down(vreg_43_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_10), .sw(sw));
	wire signed[17:0] vwire_43_11;
	reg signed[17:0] vreg_43_11;
	node n43_11(.left(vreg_42_11), .right(vreg_44_11), .up(vreg_43_12), .down(vreg_43_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_11), .sw(sw));
	wire signed[17:0] vwire_43_12;
	reg signed[17:0] vreg_43_12;
	node n43_12(.left(vreg_42_12), .right(vreg_44_12), .up(vreg_43_13), .down(vreg_43_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_12), .sw(sw));
	wire signed[17:0] vwire_43_13;
	reg signed[17:0] vreg_43_13;
	node n43_13(.left(vreg_42_13), .right(vreg_44_13), .up(vreg_43_14), .down(vreg_43_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_13), .sw(sw));
	wire signed[17:0] vwire_43_14;
	reg signed[17:0] vreg_43_14;
	node n43_14(.left(vreg_42_14), .right(vreg_44_14), .up(vreg_43_15), .down(vreg_43_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_14), .sw(sw));
	wire signed[17:0] vwire_43_15;
	reg signed[17:0] vreg_43_15;
	node n43_15(.left(vreg_42_15), .right(vreg_44_15), .up(vreg_43_16), .down(vreg_43_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_15), .sw(sw));
	wire signed[17:0] vwire_43_16;
	reg signed[17:0] vreg_43_16;
	node n43_16(.left(vreg_42_16), .right(vreg_44_16), .up(vreg_43_17), .down(vreg_43_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_16), .sw(sw));
	wire signed[17:0] vwire_43_17;
	reg signed[17:0] vreg_43_17;
	node n43_17(.left(vreg_42_17), .right(vreg_44_17), .up(vreg_43_18), .down(vreg_43_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_17), .sw(sw));
	wire signed[17:0] vwire_43_18;
	reg signed[17:0] vreg_43_18;
	node n43_18(.left(vreg_42_18), .right(vreg_44_18), .up(vreg_43_19), .down(vreg_43_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_18), .sw(sw));
	wire signed[17:0] vwire_43_19;
	reg signed[17:0] vreg_43_19;
	node n43_19(.left(vreg_42_19), .right(vreg_44_19), .up(vreg_43_20), .down(vreg_43_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_19), .sw(sw));
	wire signed[17:0] vwire_43_20;
	reg signed[17:0] vreg_43_20;
	node n43_20(.left(vreg_42_20), .right(vreg_44_20), .up(vreg_43_21), .down(vreg_43_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_20), .sw(sw));
	wire signed[17:0] vwire_43_21;
	reg signed[17:0] vreg_43_21;
	node n43_21(.left(vreg_42_21), .right(vreg_44_21), .up(vreg_43_22), .down(vreg_43_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_21), .sw(sw));
	wire signed[17:0] vwire_43_22;
	reg signed[17:0] vreg_43_22;
	node n43_22(.left(vreg_42_22), .right(vreg_44_22), .up(vreg_43_23), .down(vreg_43_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_22), .sw(sw));
	wire signed[17:0] vwire_43_23;
	reg signed[17:0] vreg_43_23;
	node n43_23(.left(vreg_42_23), .right(vreg_44_23), .up(vreg_43_24), .down(vreg_43_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_23), .sw(sw));
	wire signed[17:0] vwire_43_24;
	reg signed[17:0] vreg_43_24;
	node n43_24(.left(vreg_42_24), .right(vreg_44_24), .up(vreg_43_25), .down(vreg_43_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_24), .sw(sw));
	wire signed[17:0] vwire_43_25;
	reg signed[17:0] vreg_43_25;
	node n43_25(.left(vreg_42_25), .right(vreg_44_25), .up(vreg_43_26), .down(vreg_43_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_25), .sw(sw));
	wire signed[17:0] vwire_43_26;
	reg signed[17:0] vreg_43_26;
	node n43_26(.left(vreg_42_26), .right(vreg_44_26), .up(vreg_43_27), .down(vreg_43_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_26), .sw(sw));
	wire signed[17:0] vwire_43_27;
	reg signed[17:0] vreg_43_27;
	node n43_27(.left(vreg_42_27), .right(vreg_44_27), .up(vreg_43_28), .down(vreg_43_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_27), .sw(sw));
	wire signed[17:0] vwire_43_28;
	reg signed[17:0] vreg_43_28;
	node n43_28(.left(vreg_42_28), .right(vreg_44_28), .up(vreg_43_29), .down(vreg_43_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_28), .sw(sw));
	wire signed[17:0] vwire_43_29;
	reg signed[17:0] vreg_43_29;
	node n43_29(.left(vreg_42_29), .right(vreg_44_29), .up(vreg_43_30), .down(vreg_43_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_29), .sw(sw));
	wire signed[17:0] vwire_43_30;
	reg signed[17:0] vreg_43_30;
	node n43_30(.left(vreg_42_30), .right(vreg_44_30), .up(vreg_43_31), .down(vreg_43_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_30), .sw(sw));
	wire signed[17:0] vwire_43_31;
	reg signed[17:0] vreg_43_31;
	node n43_31(.left(vreg_42_31), .right(vreg_44_31), .up(vreg_43_32), .down(vreg_43_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_31), .sw(sw));
	wire signed[17:0] vwire_43_32;
	reg signed[17:0] vreg_43_32;
	node n43_32(.left(vreg_42_32), .right(vreg_44_32), .up(vreg_43_33), .down(vreg_43_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_32), .sw(sw));
	wire signed[17:0] vwire_43_33;
	reg signed[17:0] vreg_43_33;
	node n43_33(.left(vreg_42_33), .right(vreg_44_33), .up(vreg_43_34), .down(vreg_43_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_33), .sw(sw));
	wire signed[17:0] vwire_43_34;
	reg signed[17:0] vreg_43_34;
	node n43_34(.left(vreg_42_34), .right(vreg_44_34), .up(vreg_43_35), .down(vreg_43_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_34), .sw(sw));
	wire signed[17:0] vwire_43_35;
	reg signed[17:0] vreg_43_35;
	node n43_35(.left(vreg_42_35), .right(vreg_44_35), .up(vreg_43_36), .down(vreg_43_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_35), .sw(sw));
	wire signed[17:0] vwire_43_36;
	reg signed[17:0] vreg_43_36;
	node n43_36(.left(vreg_42_36), .right(vreg_44_36), .up(vreg_43_37), .down(vreg_43_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_36), .sw(sw));
	wire signed[17:0] vwire_43_37;
	reg signed[17:0] vreg_43_37;
	node n43_37(.left(vreg_42_37), .right(vreg_44_37), .up(vreg_43_38), .down(vreg_43_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_37), .sw(sw));
	wire signed[17:0] vwire_43_38;
	reg signed[17:0] vreg_43_38;
	node n43_38(.left(vreg_42_38), .right(vreg_44_38), .up(vreg_43_39), .down(vreg_43_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_38), .sw(sw));
	wire signed[17:0] vwire_43_39;
	reg signed[17:0] vreg_43_39;
	node n43_39(.left(vreg_42_39), .right(vreg_44_39), .up(vreg_43_40), .down(vreg_43_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_39), .sw(sw));
	wire signed[17:0] vwire_43_40;
	reg signed[17:0] vreg_43_40;
	node n43_40(.left(vreg_42_40), .right(vreg_44_40), .up(vreg_43_41), .down(vreg_43_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_40), .sw(sw));
	wire signed[17:0] vwire_43_41;
	reg signed[17:0] vreg_43_41;
	node n43_41(.left(vreg_42_41), .right(vreg_44_41), .up(vreg_43_42), .down(vreg_43_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_41), .sw(sw));
	wire signed[17:0] vwire_43_42;
	reg signed[17:0] vreg_43_42;
	node n43_42(.left(vreg_42_42), .right(vreg_44_42), .up(vreg_43_43), .down(vreg_43_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_42), .sw(sw));
	wire signed[17:0] vwire_43_43;
	reg signed[17:0] vreg_43_43;
	node n43_43(.left(vreg_42_43), .right(vreg_44_43), .up(vreg_43_44), .down(vreg_43_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_43), .sw(sw));
	wire signed[17:0] vwire_43_44;
	reg signed[17:0] vreg_43_44;
	node n43_44(.left(vreg_42_44), .right(vreg_44_44), .up(vreg_43_45), .down(vreg_43_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_44), .sw(sw));
	wire signed[17:0] vwire_43_45;
	reg signed[17:0] vreg_43_45;
	node n43_45(.left(vreg_42_45), .right(vreg_44_45), .up(vreg_43_46), .down(vreg_43_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_45), .sw(sw));
	wire signed[17:0] vwire_43_46;
	reg signed[17:0] vreg_43_46;
	node n43_46(.left(vreg_42_46), .right(vreg_44_46), .up(vreg_43_47), .down(vreg_43_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_46), .sw(sw));
	wire signed[17:0] vwire_43_47;
	reg signed[17:0] vreg_43_47;
	node n43_47(.left(vreg_42_47), .right(vreg_44_47), .up(vreg_43_48), .down(vreg_43_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_47), .sw(sw));
	wire signed[17:0] vwire_43_48;
	reg signed[17:0] vreg_43_48;
	node n43_48(.left(vreg_42_48), .right(vreg_44_48), .up(vreg_43_49), .down(vreg_43_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_48), .sw(sw));
	wire signed[17:0] vwire_43_49;
	reg signed[17:0] vreg_43_49;
	node n43_49(.left(vreg_42_49), .right(vreg_44_49), .up(18'b0), .down(vreg_43_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_43_49), .sw(sw));
	wire signed[17:0] vwire_44_0;
	reg signed[17:0] vreg_44_0;
	node n44_0(.left(vreg_43_0), .right(vreg_45_0), .up(vreg_44_1), .down(vreg_44_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_0), .sw(sw));
	wire signed[17:0] vwire_44_1;
	reg signed[17:0] vreg_44_1;
	node n44_1(.left(vreg_43_1), .right(vreg_45_1), .up(vreg_44_2), .down(vreg_44_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_1), .sw(sw));
	wire signed[17:0] vwire_44_2;
	reg signed[17:0] vreg_44_2;
	node n44_2(.left(vreg_43_2), .right(vreg_45_2), .up(vreg_44_3), .down(vreg_44_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_2), .sw(sw));
	wire signed[17:0] vwire_44_3;
	reg signed[17:0] vreg_44_3;
	node n44_3(.left(vreg_43_3), .right(vreg_45_3), .up(vreg_44_4), .down(vreg_44_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_3), .sw(sw));
	wire signed[17:0] vwire_44_4;
	reg signed[17:0] vreg_44_4;
	node n44_4(.left(vreg_43_4), .right(vreg_45_4), .up(vreg_44_5), .down(vreg_44_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_4), .sw(sw));
	wire signed[17:0] vwire_44_5;
	reg signed[17:0] vreg_44_5;
	node n44_5(.left(vreg_43_5), .right(vreg_45_5), .up(vreg_44_6), .down(vreg_44_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_5), .sw(sw));
	wire signed[17:0] vwire_44_6;
	reg signed[17:0] vreg_44_6;
	node n44_6(.left(vreg_43_6), .right(vreg_45_6), .up(vreg_44_7), .down(vreg_44_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_6), .sw(sw));
	wire signed[17:0] vwire_44_7;
	reg signed[17:0] vreg_44_7;
	node n44_7(.left(vreg_43_7), .right(vreg_45_7), .up(vreg_44_8), .down(vreg_44_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_7), .sw(sw));
	wire signed[17:0] vwire_44_8;
	reg signed[17:0] vreg_44_8;
	node n44_8(.left(vreg_43_8), .right(vreg_45_8), .up(vreg_44_9), .down(vreg_44_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_8), .sw(sw));
	wire signed[17:0] vwire_44_9;
	reg signed[17:0] vreg_44_9;
	node n44_9(.left(vreg_43_9), .right(vreg_45_9), .up(vreg_44_10), .down(vreg_44_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_9), .sw(sw));
	wire signed[17:0] vwire_44_10;
	reg signed[17:0] vreg_44_10;
	node n44_10(.left(vreg_43_10), .right(vreg_45_10), .up(vreg_44_11), .down(vreg_44_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_10), .sw(sw));
	wire signed[17:0] vwire_44_11;
	reg signed[17:0] vreg_44_11;
	node n44_11(.left(vreg_43_11), .right(vreg_45_11), .up(vreg_44_12), .down(vreg_44_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_11), .sw(sw));
	wire signed[17:0] vwire_44_12;
	reg signed[17:0] vreg_44_12;
	node n44_12(.left(vreg_43_12), .right(vreg_45_12), .up(vreg_44_13), .down(vreg_44_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_12), .sw(sw));
	wire signed[17:0] vwire_44_13;
	reg signed[17:0] vreg_44_13;
	node n44_13(.left(vreg_43_13), .right(vreg_45_13), .up(vreg_44_14), .down(vreg_44_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_13), .sw(sw));
	wire signed[17:0] vwire_44_14;
	reg signed[17:0] vreg_44_14;
	node n44_14(.left(vreg_43_14), .right(vreg_45_14), .up(vreg_44_15), .down(vreg_44_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_14), .sw(sw));
	wire signed[17:0] vwire_44_15;
	reg signed[17:0] vreg_44_15;
	node n44_15(.left(vreg_43_15), .right(vreg_45_15), .up(vreg_44_16), .down(vreg_44_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_15), .sw(sw));
	wire signed[17:0] vwire_44_16;
	reg signed[17:0] vreg_44_16;
	node n44_16(.left(vreg_43_16), .right(vreg_45_16), .up(vreg_44_17), .down(vreg_44_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_16), .sw(sw));
	wire signed[17:0] vwire_44_17;
	reg signed[17:0] vreg_44_17;
	node n44_17(.left(vreg_43_17), .right(vreg_45_17), .up(vreg_44_18), .down(vreg_44_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_17), .sw(sw));
	wire signed[17:0] vwire_44_18;
	reg signed[17:0] vreg_44_18;
	node n44_18(.left(vreg_43_18), .right(vreg_45_18), .up(vreg_44_19), .down(vreg_44_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_18), .sw(sw));
	wire signed[17:0] vwire_44_19;
	reg signed[17:0] vreg_44_19;
	node n44_19(.left(vreg_43_19), .right(vreg_45_19), .up(vreg_44_20), .down(vreg_44_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_19), .sw(sw));
	wire signed[17:0] vwire_44_20;
	reg signed[17:0] vreg_44_20;
	node n44_20(.left(vreg_43_20), .right(vreg_45_20), .up(vreg_44_21), .down(vreg_44_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_20), .sw(sw));
	wire signed[17:0] vwire_44_21;
	reg signed[17:0] vreg_44_21;
	node n44_21(.left(vreg_43_21), .right(vreg_45_21), .up(vreg_44_22), .down(vreg_44_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_21), .sw(sw));
	wire signed[17:0] vwire_44_22;
	reg signed[17:0] vreg_44_22;
	node n44_22(.left(vreg_43_22), .right(vreg_45_22), .up(vreg_44_23), .down(vreg_44_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_22), .sw(sw));
	wire signed[17:0] vwire_44_23;
	reg signed[17:0] vreg_44_23;
	node n44_23(.left(vreg_43_23), .right(vreg_45_23), .up(vreg_44_24), .down(vreg_44_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_23), .sw(sw));
	wire signed[17:0] vwire_44_24;
	reg signed[17:0] vreg_44_24;
	node n44_24(.left(vreg_43_24), .right(vreg_45_24), .up(vreg_44_25), .down(vreg_44_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_24), .sw(sw));
	wire signed[17:0] vwire_44_25;
	reg signed[17:0] vreg_44_25;
	node n44_25(.left(vreg_43_25), .right(vreg_45_25), .up(vreg_44_26), .down(vreg_44_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_25), .sw(sw));
	wire signed[17:0] vwire_44_26;
	reg signed[17:0] vreg_44_26;
	node n44_26(.left(vreg_43_26), .right(vreg_45_26), .up(vreg_44_27), .down(vreg_44_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_26), .sw(sw));
	wire signed[17:0] vwire_44_27;
	reg signed[17:0] vreg_44_27;
	node n44_27(.left(vreg_43_27), .right(vreg_45_27), .up(vreg_44_28), .down(vreg_44_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_27), .sw(sw));
	wire signed[17:0] vwire_44_28;
	reg signed[17:0] vreg_44_28;
	node n44_28(.left(vreg_43_28), .right(vreg_45_28), .up(vreg_44_29), .down(vreg_44_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_28), .sw(sw));
	wire signed[17:0] vwire_44_29;
	reg signed[17:0] vreg_44_29;
	node n44_29(.left(vreg_43_29), .right(vreg_45_29), .up(vreg_44_30), .down(vreg_44_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_29), .sw(sw));
	wire signed[17:0] vwire_44_30;
	reg signed[17:0] vreg_44_30;
	node n44_30(.left(vreg_43_30), .right(vreg_45_30), .up(vreg_44_31), .down(vreg_44_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_30), .sw(sw));
	wire signed[17:0] vwire_44_31;
	reg signed[17:0] vreg_44_31;
	node n44_31(.left(vreg_43_31), .right(vreg_45_31), .up(vreg_44_32), .down(vreg_44_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_31), .sw(sw));
	wire signed[17:0] vwire_44_32;
	reg signed[17:0] vreg_44_32;
	node n44_32(.left(vreg_43_32), .right(vreg_45_32), .up(vreg_44_33), .down(vreg_44_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_32), .sw(sw));
	wire signed[17:0] vwire_44_33;
	reg signed[17:0] vreg_44_33;
	node n44_33(.left(vreg_43_33), .right(vreg_45_33), .up(vreg_44_34), .down(vreg_44_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_33), .sw(sw));
	wire signed[17:0] vwire_44_34;
	reg signed[17:0] vreg_44_34;
	node n44_34(.left(vreg_43_34), .right(vreg_45_34), .up(vreg_44_35), .down(vreg_44_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_34), .sw(sw));
	wire signed[17:0] vwire_44_35;
	reg signed[17:0] vreg_44_35;
	node n44_35(.left(vreg_43_35), .right(vreg_45_35), .up(vreg_44_36), .down(vreg_44_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_35), .sw(sw));
	wire signed[17:0] vwire_44_36;
	reg signed[17:0] vreg_44_36;
	node n44_36(.left(vreg_43_36), .right(vreg_45_36), .up(vreg_44_37), .down(vreg_44_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_36), .sw(sw));
	wire signed[17:0] vwire_44_37;
	reg signed[17:0] vreg_44_37;
	node n44_37(.left(vreg_43_37), .right(vreg_45_37), .up(vreg_44_38), .down(vreg_44_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_37), .sw(sw));
	wire signed[17:0] vwire_44_38;
	reg signed[17:0] vreg_44_38;
	node n44_38(.left(vreg_43_38), .right(vreg_45_38), .up(vreg_44_39), .down(vreg_44_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_38), .sw(sw));
	wire signed[17:0] vwire_44_39;
	reg signed[17:0] vreg_44_39;
	node n44_39(.left(vreg_43_39), .right(vreg_45_39), .up(vreg_44_40), .down(vreg_44_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_39), .sw(sw));
	wire signed[17:0] vwire_44_40;
	reg signed[17:0] vreg_44_40;
	node n44_40(.left(vreg_43_40), .right(vreg_45_40), .up(vreg_44_41), .down(vreg_44_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_40), .sw(sw));
	wire signed[17:0] vwire_44_41;
	reg signed[17:0] vreg_44_41;
	node n44_41(.left(vreg_43_41), .right(vreg_45_41), .up(vreg_44_42), .down(vreg_44_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_41), .sw(sw));
	wire signed[17:0] vwire_44_42;
	reg signed[17:0] vreg_44_42;
	node n44_42(.left(vreg_43_42), .right(vreg_45_42), .up(vreg_44_43), .down(vreg_44_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_42), .sw(sw));
	wire signed[17:0] vwire_44_43;
	reg signed[17:0] vreg_44_43;
	node n44_43(.left(vreg_43_43), .right(vreg_45_43), .up(vreg_44_44), .down(vreg_44_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_43), .sw(sw));
	wire signed[17:0] vwire_44_44;
	reg signed[17:0] vreg_44_44;
	node n44_44(.left(vreg_43_44), .right(vreg_45_44), .up(vreg_44_45), .down(vreg_44_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_44), .sw(sw));
	wire signed[17:0] vwire_44_45;
	reg signed[17:0] vreg_44_45;
	node n44_45(.left(vreg_43_45), .right(vreg_45_45), .up(vreg_44_46), .down(vreg_44_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_45), .sw(sw));
	wire signed[17:0] vwire_44_46;
	reg signed[17:0] vreg_44_46;
	node n44_46(.left(vreg_43_46), .right(vreg_45_46), .up(vreg_44_47), .down(vreg_44_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_46), .sw(sw));
	wire signed[17:0] vwire_44_47;
	reg signed[17:0] vreg_44_47;
	node n44_47(.left(vreg_43_47), .right(vreg_45_47), .up(vreg_44_48), .down(vreg_44_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_47), .sw(sw));
	wire signed[17:0] vwire_44_48;
	reg signed[17:0] vreg_44_48;
	node n44_48(.left(vreg_43_48), .right(vreg_45_48), .up(vreg_44_49), .down(vreg_44_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_48), .sw(sw));
	wire signed[17:0] vwire_44_49;
	reg signed[17:0] vreg_44_49;
	node n44_49(.left(vreg_43_49), .right(vreg_45_49), .up(18'b0), .down(vreg_44_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_44_49), .sw(sw));
	wire signed[17:0] vwire_45_0;
	reg signed[17:0] vreg_45_0;
	node n45_0(.left(vreg_44_0), .right(vreg_46_0), .up(vreg_45_1), .down(vreg_45_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_0), .sw(sw));
	wire signed[17:0] vwire_45_1;
	reg signed[17:0] vreg_45_1;
	node n45_1(.left(vreg_44_1), .right(vreg_46_1), .up(vreg_45_2), .down(vreg_45_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_1), .sw(sw));
	wire signed[17:0] vwire_45_2;
	reg signed[17:0] vreg_45_2;
	node n45_2(.left(vreg_44_2), .right(vreg_46_2), .up(vreg_45_3), .down(vreg_45_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_2), .sw(sw));
	wire signed[17:0] vwire_45_3;
	reg signed[17:0] vreg_45_3;
	node n45_3(.left(vreg_44_3), .right(vreg_46_3), .up(vreg_45_4), .down(vreg_45_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_3), .sw(sw));
	wire signed[17:0] vwire_45_4;
	reg signed[17:0] vreg_45_4;
	node n45_4(.left(vreg_44_4), .right(vreg_46_4), .up(vreg_45_5), .down(vreg_45_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_4), .sw(sw));
	wire signed[17:0] vwire_45_5;
	reg signed[17:0] vreg_45_5;
	node n45_5(.left(vreg_44_5), .right(vreg_46_5), .up(vreg_45_6), .down(vreg_45_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_5), .sw(sw));
	wire signed[17:0] vwire_45_6;
	reg signed[17:0] vreg_45_6;
	node n45_6(.left(vreg_44_6), .right(vreg_46_6), .up(vreg_45_7), .down(vreg_45_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_6), .sw(sw));
	wire signed[17:0] vwire_45_7;
	reg signed[17:0] vreg_45_7;
	node n45_7(.left(vreg_44_7), .right(vreg_46_7), .up(vreg_45_8), .down(vreg_45_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_7), .sw(sw));
	wire signed[17:0] vwire_45_8;
	reg signed[17:0] vreg_45_8;
	node n45_8(.left(vreg_44_8), .right(vreg_46_8), .up(vreg_45_9), .down(vreg_45_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_8), .sw(sw));
	wire signed[17:0] vwire_45_9;
	reg signed[17:0] vreg_45_9;
	node n45_9(.left(vreg_44_9), .right(vreg_46_9), .up(vreg_45_10), .down(vreg_45_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_9), .sw(sw));
	wire signed[17:0] vwire_45_10;
	reg signed[17:0] vreg_45_10;
	node n45_10(.left(vreg_44_10), .right(vreg_46_10), .up(vreg_45_11), .down(vreg_45_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_10), .sw(sw));
	wire signed[17:0] vwire_45_11;
	reg signed[17:0] vreg_45_11;
	node n45_11(.left(vreg_44_11), .right(vreg_46_11), .up(vreg_45_12), .down(vreg_45_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_11), .sw(sw));
	wire signed[17:0] vwire_45_12;
	reg signed[17:0] vreg_45_12;
	node n45_12(.left(vreg_44_12), .right(vreg_46_12), .up(vreg_45_13), .down(vreg_45_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_12), .sw(sw));
	wire signed[17:0] vwire_45_13;
	reg signed[17:0] vreg_45_13;
	node n45_13(.left(vreg_44_13), .right(vreg_46_13), .up(vreg_45_14), .down(vreg_45_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_13), .sw(sw));
	wire signed[17:0] vwire_45_14;
	reg signed[17:0] vreg_45_14;
	node n45_14(.left(vreg_44_14), .right(vreg_46_14), .up(vreg_45_15), .down(vreg_45_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_14), .sw(sw));
	wire signed[17:0] vwire_45_15;
	reg signed[17:0] vreg_45_15;
	node n45_15(.left(vreg_44_15), .right(vreg_46_15), .up(vreg_45_16), .down(vreg_45_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_15), .sw(sw));
	wire signed[17:0] vwire_45_16;
	reg signed[17:0] vreg_45_16;
	node n45_16(.left(vreg_44_16), .right(vreg_46_16), .up(vreg_45_17), .down(vreg_45_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_16), .sw(sw));
	wire signed[17:0] vwire_45_17;
	reg signed[17:0] vreg_45_17;
	node n45_17(.left(vreg_44_17), .right(vreg_46_17), .up(vreg_45_18), .down(vreg_45_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_17), .sw(sw));
	wire signed[17:0] vwire_45_18;
	reg signed[17:0] vreg_45_18;
	node n45_18(.left(vreg_44_18), .right(vreg_46_18), .up(vreg_45_19), .down(vreg_45_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_18), .sw(sw));
	wire signed[17:0] vwire_45_19;
	reg signed[17:0] vreg_45_19;
	node n45_19(.left(vreg_44_19), .right(vreg_46_19), .up(vreg_45_20), .down(vreg_45_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_19), .sw(sw));
	wire signed[17:0] vwire_45_20;
	reg signed[17:0] vreg_45_20;
	node n45_20(.left(vreg_44_20), .right(vreg_46_20), .up(vreg_45_21), .down(vreg_45_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_20), .sw(sw));
	wire signed[17:0] vwire_45_21;
	reg signed[17:0] vreg_45_21;
	node n45_21(.left(vreg_44_21), .right(vreg_46_21), .up(vreg_45_22), .down(vreg_45_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_21), .sw(sw));
	wire signed[17:0] vwire_45_22;
	reg signed[17:0] vreg_45_22;
	node n45_22(.left(vreg_44_22), .right(vreg_46_22), .up(vreg_45_23), .down(vreg_45_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_22), .sw(sw));
	wire signed[17:0] vwire_45_23;
	reg signed[17:0] vreg_45_23;
	node n45_23(.left(vreg_44_23), .right(vreg_46_23), .up(vreg_45_24), .down(vreg_45_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_23), .sw(sw));
	wire signed[17:0] vwire_45_24;
	reg signed[17:0] vreg_45_24;
	node n45_24(.left(vreg_44_24), .right(vreg_46_24), .up(vreg_45_25), .down(vreg_45_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_24), .sw(sw));
	wire signed[17:0] vwire_45_25;
	reg signed[17:0] vreg_45_25;
	node n45_25(.left(vreg_44_25), .right(vreg_46_25), .up(vreg_45_26), .down(vreg_45_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_25), .sw(sw));
	wire signed[17:0] vwire_45_26;
	reg signed[17:0] vreg_45_26;
	node n45_26(.left(vreg_44_26), .right(vreg_46_26), .up(vreg_45_27), .down(vreg_45_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_26), .sw(sw));
	wire signed[17:0] vwire_45_27;
	reg signed[17:0] vreg_45_27;
	node n45_27(.left(vreg_44_27), .right(vreg_46_27), .up(vreg_45_28), .down(vreg_45_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_27), .sw(sw));
	wire signed[17:0] vwire_45_28;
	reg signed[17:0] vreg_45_28;
	node n45_28(.left(vreg_44_28), .right(vreg_46_28), .up(vreg_45_29), .down(vreg_45_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_28), .sw(sw));
	wire signed[17:0] vwire_45_29;
	reg signed[17:0] vreg_45_29;
	node n45_29(.left(vreg_44_29), .right(vreg_46_29), .up(vreg_45_30), .down(vreg_45_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_29), .sw(sw));
	wire signed[17:0] vwire_45_30;
	reg signed[17:0] vreg_45_30;
	node n45_30(.left(vreg_44_30), .right(vreg_46_30), .up(vreg_45_31), .down(vreg_45_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_30), .sw(sw));
	wire signed[17:0] vwire_45_31;
	reg signed[17:0] vreg_45_31;
	node n45_31(.left(vreg_44_31), .right(vreg_46_31), .up(vreg_45_32), .down(vreg_45_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_31), .sw(sw));
	wire signed[17:0] vwire_45_32;
	reg signed[17:0] vreg_45_32;
	node n45_32(.left(vreg_44_32), .right(vreg_46_32), .up(vreg_45_33), .down(vreg_45_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_32), .sw(sw));
	wire signed[17:0] vwire_45_33;
	reg signed[17:0] vreg_45_33;
	node n45_33(.left(vreg_44_33), .right(vreg_46_33), .up(vreg_45_34), .down(vreg_45_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_33), .sw(sw));
	wire signed[17:0] vwire_45_34;
	reg signed[17:0] vreg_45_34;
	node n45_34(.left(vreg_44_34), .right(vreg_46_34), .up(vreg_45_35), .down(vreg_45_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_34), .sw(sw));
	wire signed[17:0] vwire_45_35;
	reg signed[17:0] vreg_45_35;
	node n45_35(.left(vreg_44_35), .right(vreg_46_35), .up(vreg_45_36), .down(vreg_45_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_35), .sw(sw));
	wire signed[17:0] vwire_45_36;
	reg signed[17:0] vreg_45_36;
	node n45_36(.left(vreg_44_36), .right(vreg_46_36), .up(vreg_45_37), .down(vreg_45_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_36), .sw(sw));
	wire signed[17:0] vwire_45_37;
	reg signed[17:0] vreg_45_37;
	node n45_37(.left(vreg_44_37), .right(vreg_46_37), .up(vreg_45_38), .down(vreg_45_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_37), .sw(sw));
	wire signed[17:0] vwire_45_38;
	reg signed[17:0] vreg_45_38;
	node n45_38(.left(vreg_44_38), .right(vreg_46_38), .up(vreg_45_39), .down(vreg_45_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_38), .sw(sw));
	wire signed[17:0] vwire_45_39;
	reg signed[17:0] vreg_45_39;
	node n45_39(.left(vreg_44_39), .right(vreg_46_39), .up(vreg_45_40), .down(vreg_45_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_39), .sw(sw));
	wire signed[17:0] vwire_45_40;
	reg signed[17:0] vreg_45_40;
	node n45_40(.left(vreg_44_40), .right(vreg_46_40), .up(vreg_45_41), .down(vreg_45_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_40), .sw(sw));
	wire signed[17:0] vwire_45_41;
	reg signed[17:0] vreg_45_41;
	node n45_41(.left(vreg_44_41), .right(vreg_46_41), .up(vreg_45_42), .down(vreg_45_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_41), .sw(sw));
	wire signed[17:0] vwire_45_42;
	reg signed[17:0] vreg_45_42;
	node n45_42(.left(vreg_44_42), .right(vreg_46_42), .up(vreg_45_43), .down(vreg_45_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_42), .sw(sw));
	wire signed[17:0] vwire_45_43;
	reg signed[17:0] vreg_45_43;
	node n45_43(.left(vreg_44_43), .right(vreg_46_43), .up(vreg_45_44), .down(vreg_45_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_43), .sw(sw));
	wire signed[17:0] vwire_45_44;
	reg signed[17:0] vreg_45_44;
	node n45_44(.left(vreg_44_44), .right(vreg_46_44), .up(vreg_45_45), .down(vreg_45_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_44), .sw(sw));
	wire signed[17:0] vwire_45_45;
	reg signed[17:0] vreg_45_45;
	node n45_45(.left(vreg_44_45), .right(vreg_46_45), .up(vreg_45_46), .down(vreg_45_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_45), .sw(sw));
	wire signed[17:0] vwire_45_46;
	reg signed[17:0] vreg_45_46;
	node n45_46(.left(vreg_44_46), .right(vreg_46_46), .up(vreg_45_47), .down(vreg_45_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_46), .sw(sw));
	wire signed[17:0] vwire_45_47;
	reg signed[17:0] vreg_45_47;
	node n45_47(.left(vreg_44_47), .right(vreg_46_47), .up(vreg_45_48), .down(vreg_45_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_47), .sw(sw));
	wire signed[17:0] vwire_45_48;
	reg signed[17:0] vreg_45_48;
	node n45_48(.left(vreg_44_48), .right(vreg_46_48), .up(vreg_45_49), .down(vreg_45_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_48), .sw(sw));
	wire signed[17:0] vwire_45_49;
	reg signed[17:0] vreg_45_49;
	node n45_49(.left(vreg_44_49), .right(vreg_46_49), .up(18'b0), .down(vreg_45_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_45_49), .sw(sw));
	wire signed[17:0] vwire_46_0;
	reg signed[17:0] vreg_46_0;
	node n46_0(.left(vreg_45_0), .right(vreg_47_0), .up(vreg_46_1), .down(vreg_46_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_0), .sw(sw));
	wire signed[17:0] vwire_46_1;
	reg signed[17:0] vreg_46_1;
	node n46_1(.left(vreg_45_1), .right(vreg_47_1), .up(vreg_46_2), .down(vreg_46_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_1), .sw(sw));
	wire signed[17:0] vwire_46_2;
	reg signed[17:0] vreg_46_2;
	node n46_2(.left(vreg_45_2), .right(vreg_47_2), .up(vreg_46_3), .down(vreg_46_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_2), .sw(sw));
	wire signed[17:0] vwire_46_3;
	reg signed[17:0] vreg_46_3;
	node n46_3(.left(vreg_45_3), .right(vreg_47_3), .up(vreg_46_4), .down(vreg_46_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_3), .sw(sw));
	wire signed[17:0] vwire_46_4;
	reg signed[17:0] vreg_46_4;
	node n46_4(.left(vreg_45_4), .right(vreg_47_4), .up(vreg_46_5), .down(vreg_46_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_4), .sw(sw));
	wire signed[17:0] vwire_46_5;
	reg signed[17:0] vreg_46_5;
	node n46_5(.left(vreg_45_5), .right(vreg_47_5), .up(vreg_46_6), .down(vreg_46_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_5), .sw(sw));
	wire signed[17:0] vwire_46_6;
	reg signed[17:0] vreg_46_6;
	node n46_6(.left(vreg_45_6), .right(vreg_47_6), .up(vreg_46_7), .down(vreg_46_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_6), .sw(sw));
	wire signed[17:0] vwire_46_7;
	reg signed[17:0] vreg_46_7;
	node n46_7(.left(vreg_45_7), .right(vreg_47_7), .up(vreg_46_8), .down(vreg_46_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_7), .sw(sw));
	wire signed[17:0] vwire_46_8;
	reg signed[17:0] vreg_46_8;
	node n46_8(.left(vreg_45_8), .right(vreg_47_8), .up(vreg_46_9), .down(vreg_46_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_8), .sw(sw));
	wire signed[17:0] vwire_46_9;
	reg signed[17:0] vreg_46_9;
	node n46_9(.left(vreg_45_9), .right(vreg_47_9), .up(vreg_46_10), .down(vreg_46_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_9), .sw(sw));
	wire signed[17:0] vwire_46_10;
	reg signed[17:0] vreg_46_10;
	node n46_10(.left(vreg_45_10), .right(vreg_47_10), .up(vreg_46_11), .down(vreg_46_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_10), .sw(sw));
	wire signed[17:0] vwire_46_11;
	reg signed[17:0] vreg_46_11;
	node n46_11(.left(vreg_45_11), .right(vreg_47_11), .up(vreg_46_12), .down(vreg_46_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_11), .sw(sw));
	wire signed[17:0] vwire_46_12;
	reg signed[17:0] vreg_46_12;
	node n46_12(.left(vreg_45_12), .right(vreg_47_12), .up(vreg_46_13), .down(vreg_46_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_12), .sw(sw));
	wire signed[17:0] vwire_46_13;
	reg signed[17:0] vreg_46_13;
	node n46_13(.left(vreg_45_13), .right(vreg_47_13), .up(vreg_46_14), .down(vreg_46_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_13), .sw(sw));
	wire signed[17:0] vwire_46_14;
	reg signed[17:0] vreg_46_14;
	node n46_14(.left(vreg_45_14), .right(vreg_47_14), .up(vreg_46_15), .down(vreg_46_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_14), .sw(sw));
	wire signed[17:0] vwire_46_15;
	reg signed[17:0] vreg_46_15;
	node n46_15(.left(vreg_45_15), .right(vreg_47_15), .up(vreg_46_16), .down(vreg_46_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_15), .sw(sw));
	wire signed[17:0] vwire_46_16;
	reg signed[17:0] vreg_46_16;
	node n46_16(.left(vreg_45_16), .right(vreg_47_16), .up(vreg_46_17), .down(vreg_46_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_16), .sw(sw));
	wire signed[17:0] vwire_46_17;
	reg signed[17:0] vreg_46_17;
	node n46_17(.left(vreg_45_17), .right(vreg_47_17), .up(vreg_46_18), .down(vreg_46_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_17), .sw(sw));
	wire signed[17:0] vwire_46_18;
	reg signed[17:0] vreg_46_18;
	node n46_18(.left(vreg_45_18), .right(vreg_47_18), .up(vreg_46_19), .down(vreg_46_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_18), .sw(sw));
	wire signed[17:0] vwire_46_19;
	reg signed[17:0] vreg_46_19;
	node n46_19(.left(vreg_45_19), .right(vreg_47_19), .up(vreg_46_20), .down(vreg_46_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_19), .sw(sw));
	wire signed[17:0] vwire_46_20;
	reg signed[17:0] vreg_46_20;
	node n46_20(.left(vreg_45_20), .right(vreg_47_20), .up(vreg_46_21), .down(vreg_46_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_20), .sw(sw));
	wire signed[17:0] vwire_46_21;
	reg signed[17:0] vreg_46_21;
	node n46_21(.left(vreg_45_21), .right(vreg_47_21), .up(vreg_46_22), .down(vreg_46_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_21), .sw(sw));
	wire signed[17:0] vwire_46_22;
	reg signed[17:0] vreg_46_22;
	node n46_22(.left(vreg_45_22), .right(vreg_47_22), .up(vreg_46_23), .down(vreg_46_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_22), .sw(sw));
	wire signed[17:0] vwire_46_23;
	reg signed[17:0] vreg_46_23;
	node n46_23(.left(vreg_45_23), .right(vreg_47_23), .up(vreg_46_24), .down(vreg_46_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_23), .sw(sw));
	wire signed[17:0] vwire_46_24;
	reg signed[17:0] vreg_46_24;
	node n46_24(.left(vreg_45_24), .right(vreg_47_24), .up(vreg_46_25), .down(vreg_46_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_24), .sw(sw));
	wire signed[17:0] vwire_46_25;
	reg signed[17:0] vreg_46_25;
	node n46_25(.left(vreg_45_25), .right(vreg_47_25), .up(vreg_46_26), .down(vreg_46_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_25), .sw(sw));
	wire signed[17:0] vwire_46_26;
	reg signed[17:0] vreg_46_26;
	node n46_26(.left(vreg_45_26), .right(vreg_47_26), .up(vreg_46_27), .down(vreg_46_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_26), .sw(sw));
	wire signed[17:0] vwire_46_27;
	reg signed[17:0] vreg_46_27;
	node n46_27(.left(vreg_45_27), .right(vreg_47_27), .up(vreg_46_28), .down(vreg_46_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_27), .sw(sw));
	wire signed[17:0] vwire_46_28;
	reg signed[17:0] vreg_46_28;
	node n46_28(.left(vreg_45_28), .right(vreg_47_28), .up(vreg_46_29), .down(vreg_46_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_28), .sw(sw));
	wire signed[17:0] vwire_46_29;
	reg signed[17:0] vreg_46_29;
	node n46_29(.left(vreg_45_29), .right(vreg_47_29), .up(vreg_46_30), .down(vreg_46_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_29), .sw(sw));
	wire signed[17:0] vwire_46_30;
	reg signed[17:0] vreg_46_30;
	node n46_30(.left(vreg_45_30), .right(vreg_47_30), .up(vreg_46_31), .down(vreg_46_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_30), .sw(sw));
	wire signed[17:0] vwire_46_31;
	reg signed[17:0] vreg_46_31;
	node n46_31(.left(vreg_45_31), .right(vreg_47_31), .up(vreg_46_32), .down(vreg_46_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_31), .sw(sw));
	wire signed[17:0] vwire_46_32;
	reg signed[17:0] vreg_46_32;
	node n46_32(.left(vreg_45_32), .right(vreg_47_32), .up(vreg_46_33), .down(vreg_46_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_32), .sw(sw));
	wire signed[17:0] vwire_46_33;
	reg signed[17:0] vreg_46_33;
	node n46_33(.left(vreg_45_33), .right(vreg_47_33), .up(vreg_46_34), .down(vreg_46_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_33), .sw(sw));
	wire signed[17:0] vwire_46_34;
	reg signed[17:0] vreg_46_34;
	node n46_34(.left(vreg_45_34), .right(vreg_47_34), .up(vreg_46_35), .down(vreg_46_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_34), .sw(sw));
	wire signed[17:0] vwire_46_35;
	reg signed[17:0] vreg_46_35;
	node n46_35(.left(vreg_45_35), .right(vreg_47_35), .up(vreg_46_36), .down(vreg_46_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_35), .sw(sw));
	wire signed[17:0] vwire_46_36;
	reg signed[17:0] vreg_46_36;
	node n46_36(.left(vreg_45_36), .right(vreg_47_36), .up(vreg_46_37), .down(vreg_46_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_36), .sw(sw));
	wire signed[17:0] vwire_46_37;
	reg signed[17:0] vreg_46_37;
	node n46_37(.left(vreg_45_37), .right(vreg_47_37), .up(vreg_46_38), .down(vreg_46_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_37), .sw(sw));
	wire signed[17:0] vwire_46_38;
	reg signed[17:0] vreg_46_38;
	node n46_38(.left(vreg_45_38), .right(vreg_47_38), .up(vreg_46_39), .down(vreg_46_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_38), .sw(sw));
	wire signed[17:0] vwire_46_39;
	reg signed[17:0] vreg_46_39;
	node n46_39(.left(vreg_45_39), .right(vreg_47_39), .up(vreg_46_40), .down(vreg_46_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_39), .sw(sw));
	wire signed[17:0] vwire_46_40;
	reg signed[17:0] vreg_46_40;
	node n46_40(.left(vreg_45_40), .right(vreg_47_40), .up(vreg_46_41), .down(vreg_46_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_40), .sw(sw));
	wire signed[17:0] vwire_46_41;
	reg signed[17:0] vreg_46_41;
	node n46_41(.left(vreg_45_41), .right(vreg_47_41), .up(vreg_46_42), .down(vreg_46_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_41), .sw(sw));
	wire signed[17:0] vwire_46_42;
	reg signed[17:0] vreg_46_42;
	node n46_42(.left(vreg_45_42), .right(vreg_47_42), .up(vreg_46_43), .down(vreg_46_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_42), .sw(sw));
	wire signed[17:0] vwire_46_43;
	reg signed[17:0] vreg_46_43;
	node n46_43(.left(vreg_45_43), .right(vreg_47_43), .up(vreg_46_44), .down(vreg_46_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_43), .sw(sw));
	wire signed[17:0] vwire_46_44;
	reg signed[17:0] vreg_46_44;
	node n46_44(.left(vreg_45_44), .right(vreg_47_44), .up(vreg_46_45), .down(vreg_46_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_44), .sw(sw));
	wire signed[17:0] vwire_46_45;
	reg signed[17:0] vreg_46_45;
	node n46_45(.left(vreg_45_45), .right(vreg_47_45), .up(vreg_46_46), .down(vreg_46_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_45), .sw(sw));
	wire signed[17:0] vwire_46_46;
	reg signed[17:0] vreg_46_46;
	node n46_46(.left(vreg_45_46), .right(vreg_47_46), .up(vreg_46_47), .down(vreg_46_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_46), .sw(sw));
	wire signed[17:0] vwire_46_47;
	reg signed[17:0] vreg_46_47;
	node n46_47(.left(vreg_45_47), .right(vreg_47_47), .up(vreg_46_48), .down(vreg_46_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_47), .sw(sw));
	wire signed[17:0] vwire_46_48;
	reg signed[17:0] vreg_46_48;
	node n46_48(.left(vreg_45_48), .right(vreg_47_48), .up(vreg_46_49), .down(vreg_46_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_48), .sw(sw));
	wire signed[17:0] vwire_46_49;
	reg signed[17:0] vreg_46_49;
	node n46_49(.left(vreg_45_49), .right(vreg_47_49), .up(18'b0), .down(vreg_46_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_46_49), .sw(sw));
	wire signed[17:0] vwire_47_0;
	reg signed[17:0] vreg_47_0;
	node n47_0(.left(vreg_46_0), .right(vreg_48_0), .up(vreg_47_1), .down(vreg_47_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_0), .sw(sw));
	wire signed[17:0] vwire_47_1;
	reg signed[17:0] vreg_47_1;
	node n47_1(.left(vreg_46_1), .right(vreg_48_1), .up(vreg_47_2), .down(vreg_47_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_1), .sw(sw));
	wire signed[17:0] vwire_47_2;
	reg signed[17:0] vreg_47_2;
	node n47_2(.left(vreg_46_2), .right(vreg_48_2), .up(vreg_47_3), .down(vreg_47_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_2), .sw(sw));
	wire signed[17:0] vwire_47_3;
	reg signed[17:0] vreg_47_3;
	node n47_3(.left(vreg_46_3), .right(vreg_48_3), .up(vreg_47_4), .down(vreg_47_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_3), .sw(sw));
	wire signed[17:0] vwire_47_4;
	reg signed[17:0] vreg_47_4;
	node n47_4(.left(vreg_46_4), .right(vreg_48_4), .up(vreg_47_5), .down(vreg_47_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_4), .sw(sw));
	wire signed[17:0] vwire_47_5;
	reg signed[17:0] vreg_47_5;
	node n47_5(.left(vreg_46_5), .right(vreg_48_5), .up(vreg_47_6), .down(vreg_47_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_5), .sw(sw));
	wire signed[17:0] vwire_47_6;
	reg signed[17:0] vreg_47_6;
	node n47_6(.left(vreg_46_6), .right(vreg_48_6), .up(vreg_47_7), .down(vreg_47_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_6), .sw(sw));
	wire signed[17:0] vwire_47_7;
	reg signed[17:0] vreg_47_7;
	node n47_7(.left(vreg_46_7), .right(vreg_48_7), .up(vreg_47_8), .down(vreg_47_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_7), .sw(sw));
	wire signed[17:0] vwire_47_8;
	reg signed[17:0] vreg_47_8;
	node n47_8(.left(vreg_46_8), .right(vreg_48_8), .up(vreg_47_9), .down(vreg_47_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_8), .sw(sw));
	wire signed[17:0] vwire_47_9;
	reg signed[17:0] vreg_47_9;
	node n47_9(.left(vreg_46_9), .right(vreg_48_9), .up(vreg_47_10), .down(vreg_47_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_9), .sw(sw));
	wire signed[17:0] vwire_47_10;
	reg signed[17:0] vreg_47_10;
	node n47_10(.left(vreg_46_10), .right(vreg_48_10), .up(vreg_47_11), .down(vreg_47_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_10), .sw(sw));
	wire signed[17:0] vwire_47_11;
	reg signed[17:0] vreg_47_11;
	node n47_11(.left(vreg_46_11), .right(vreg_48_11), .up(vreg_47_12), .down(vreg_47_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_11), .sw(sw));
	wire signed[17:0] vwire_47_12;
	reg signed[17:0] vreg_47_12;
	node n47_12(.left(vreg_46_12), .right(vreg_48_12), .up(vreg_47_13), .down(vreg_47_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_12), .sw(sw));
	wire signed[17:0] vwire_47_13;
	reg signed[17:0] vreg_47_13;
	node n47_13(.left(vreg_46_13), .right(vreg_48_13), .up(vreg_47_14), .down(vreg_47_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_13), .sw(sw));
	wire signed[17:0] vwire_47_14;
	reg signed[17:0] vreg_47_14;
	node n47_14(.left(vreg_46_14), .right(vreg_48_14), .up(vreg_47_15), .down(vreg_47_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_14), .sw(sw));
	wire signed[17:0] vwire_47_15;
	reg signed[17:0] vreg_47_15;
	node n47_15(.left(vreg_46_15), .right(vreg_48_15), .up(vreg_47_16), .down(vreg_47_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_15), .sw(sw));
	wire signed[17:0] vwire_47_16;
	reg signed[17:0] vreg_47_16;
	node n47_16(.left(vreg_46_16), .right(vreg_48_16), .up(vreg_47_17), .down(vreg_47_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_16), .sw(sw));
	wire signed[17:0] vwire_47_17;
	reg signed[17:0] vreg_47_17;
	node n47_17(.left(vreg_46_17), .right(vreg_48_17), .up(vreg_47_18), .down(vreg_47_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_17), .sw(sw));
	wire signed[17:0] vwire_47_18;
	reg signed[17:0] vreg_47_18;
	node n47_18(.left(vreg_46_18), .right(vreg_48_18), .up(vreg_47_19), .down(vreg_47_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_18), .sw(sw));
	wire signed[17:0] vwire_47_19;
	reg signed[17:0] vreg_47_19;
	node n47_19(.left(vreg_46_19), .right(vreg_48_19), .up(vreg_47_20), .down(vreg_47_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_19), .sw(sw));
	wire signed[17:0] vwire_47_20;
	reg signed[17:0] vreg_47_20;
	node n47_20(.left(vreg_46_20), .right(vreg_48_20), .up(vreg_47_21), .down(vreg_47_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_20), .sw(sw));
	wire signed[17:0] vwire_47_21;
	reg signed[17:0] vreg_47_21;
	node n47_21(.left(vreg_46_21), .right(vreg_48_21), .up(vreg_47_22), .down(vreg_47_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_21), .sw(sw));
	wire signed[17:0] vwire_47_22;
	reg signed[17:0] vreg_47_22;
	node n47_22(.left(vreg_46_22), .right(vreg_48_22), .up(vreg_47_23), .down(vreg_47_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_22), .sw(sw));
	wire signed[17:0] vwire_47_23;
	reg signed[17:0] vreg_47_23;
	node n47_23(.left(vreg_46_23), .right(vreg_48_23), .up(vreg_47_24), .down(vreg_47_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_23), .sw(sw));
	wire signed[17:0] vwire_47_24;
	reg signed[17:0] vreg_47_24;
	node n47_24(.left(vreg_46_24), .right(vreg_48_24), .up(vreg_47_25), .down(vreg_47_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_24), .sw(sw));
	wire signed[17:0] vwire_47_25;
	reg signed[17:0] vreg_47_25;
	node n47_25(.left(vreg_46_25), .right(vreg_48_25), .up(vreg_47_26), .down(vreg_47_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_25), .sw(sw));
	wire signed[17:0] vwire_47_26;
	reg signed[17:0] vreg_47_26;
	node n47_26(.left(vreg_46_26), .right(vreg_48_26), .up(vreg_47_27), .down(vreg_47_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_26), .sw(sw));
	wire signed[17:0] vwire_47_27;
	reg signed[17:0] vreg_47_27;
	node n47_27(.left(vreg_46_27), .right(vreg_48_27), .up(vreg_47_28), .down(vreg_47_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_27), .sw(sw));
	wire signed[17:0] vwire_47_28;
	reg signed[17:0] vreg_47_28;
	node n47_28(.left(vreg_46_28), .right(vreg_48_28), .up(vreg_47_29), .down(vreg_47_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_28), .sw(sw));
	wire signed[17:0] vwire_47_29;
	reg signed[17:0] vreg_47_29;
	node n47_29(.left(vreg_46_29), .right(vreg_48_29), .up(vreg_47_30), .down(vreg_47_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_29), .sw(sw));
	wire signed[17:0] vwire_47_30;
	reg signed[17:0] vreg_47_30;
	node n47_30(.left(vreg_46_30), .right(vreg_48_30), .up(vreg_47_31), .down(vreg_47_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_30), .sw(sw));
	wire signed[17:0] vwire_47_31;
	reg signed[17:0] vreg_47_31;
	node n47_31(.left(vreg_46_31), .right(vreg_48_31), .up(vreg_47_32), .down(vreg_47_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_31), .sw(sw));
	wire signed[17:0] vwire_47_32;
	reg signed[17:0] vreg_47_32;
	node n47_32(.left(vreg_46_32), .right(vreg_48_32), .up(vreg_47_33), .down(vreg_47_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_32), .sw(sw));
	wire signed[17:0] vwire_47_33;
	reg signed[17:0] vreg_47_33;
	node n47_33(.left(vreg_46_33), .right(vreg_48_33), .up(vreg_47_34), .down(vreg_47_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_33), .sw(sw));
	wire signed[17:0] vwire_47_34;
	reg signed[17:0] vreg_47_34;
	node n47_34(.left(vreg_46_34), .right(vreg_48_34), .up(vreg_47_35), .down(vreg_47_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_34), .sw(sw));
	wire signed[17:0] vwire_47_35;
	reg signed[17:0] vreg_47_35;
	node n47_35(.left(vreg_46_35), .right(vreg_48_35), .up(vreg_47_36), .down(vreg_47_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_35), .sw(sw));
	wire signed[17:0] vwire_47_36;
	reg signed[17:0] vreg_47_36;
	node n47_36(.left(vreg_46_36), .right(vreg_48_36), .up(vreg_47_37), .down(vreg_47_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_36), .sw(sw));
	wire signed[17:0] vwire_47_37;
	reg signed[17:0] vreg_47_37;
	node n47_37(.left(vreg_46_37), .right(vreg_48_37), .up(vreg_47_38), .down(vreg_47_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_37), .sw(sw));
	wire signed[17:0] vwire_47_38;
	reg signed[17:0] vreg_47_38;
	node n47_38(.left(vreg_46_38), .right(vreg_48_38), .up(vreg_47_39), .down(vreg_47_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_38), .sw(sw));
	wire signed[17:0] vwire_47_39;
	reg signed[17:0] vreg_47_39;
	node n47_39(.left(vreg_46_39), .right(vreg_48_39), .up(vreg_47_40), .down(vreg_47_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_39), .sw(sw));
	wire signed[17:0] vwire_47_40;
	reg signed[17:0] vreg_47_40;
	node n47_40(.left(vreg_46_40), .right(vreg_48_40), .up(vreg_47_41), .down(vreg_47_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_40), .sw(sw));
	wire signed[17:0] vwire_47_41;
	reg signed[17:0] vreg_47_41;
	node n47_41(.left(vreg_46_41), .right(vreg_48_41), .up(vreg_47_42), .down(vreg_47_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_41), .sw(sw));
	wire signed[17:0] vwire_47_42;
	reg signed[17:0] vreg_47_42;
	node n47_42(.left(vreg_46_42), .right(vreg_48_42), .up(vreg_47_43), .down(vreg_47_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_42), .sw(sw));
	wire signed[17:0] vwire_47_43;
	reg signed[17:0] vreg_47_43;
	node n47_43(.left(vreg_46_43), .right(vreg_48_43), .up(vreg_47_44), .down(vreg_47_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_43), .sw(sw));
	wire signed[17:0] vwire_47_44;
	reg signed[17:0] vreg_47_44;
	node n47_44(.left(vreg_46_44), .right(vreg_48_44), .up(vreg_47_45), .down(vreg_47_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_44), .sw(sw));
	wire signed[17:0] vwire_47_45;
	reg signed[17:0] vreg_47_45;
	node n47_45(.left(vreg_46_45), .right(vreg_48_45), .up(vreg_47_46), .down(vreg_47_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_45), .sw(sw));
	wire signed[17:0] vwire_47_46;
	reg signed[17:0] vreg_47_46;
	node n47_46(.left(vreg_46_46), .right(vreg_48_46), .up(vreg_47_47), .down(vreg_47_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_46), .sw(sw));
	wire signed[17:0] vwire_47_47;
	reg signed[17:0] vreg_47_47;
	node n47_47(.left(vreg_46_47), .right(vreg_48_47), .up(vreg_47_48), .down(vreg_47_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_47), .sw(sw));
	wire signed[17:0] vwire_47_48;
	reg signed[17:0] vreg_47_48;
	node n47_48(.left(vreg_46_48), .right(vreg_48_48), .up(vreg_47_49), .down(vreg_47_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_48), .sw(sw));
	wire signed[17:0] vwire_47_49;
	reg signed[17:0] vreg_47_49;
	node n47_49(.left(vreg_46_49), .right(vreg_48_49), .up(18'b0), .down(vreg_47_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_47_49), .sw(sw));
	wire signed[17:0] vwire_48_0;
	reg signed[17:0] vreg_48_0;
	node n48_0(.left(vreg_47_0), .right(vreg_49_0), .up(vreg_48_1), .down(vreg_48_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_0), .sw(sw));
	wire signed[17:0] vwire_48_1;
	reg signed[17:0] vreg_48_1;
	node n48_1(.left(vreg_47_1), .right(vreg_49_1), .up(vreg_48_2), .down(vreg_48_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_1), .sw(sw));
	wire signed[17:0] vwire_48_2;
	reg signed[17:0] vreg_48_2;
	node n48_2(.left(vreg_47_2), .right(vreg_49_2), .up(vreg_48_3), .down(vreg_48_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_2), .sw(sw));
	wire signed[17:0] vwire_48_3;
	reg signed[17:0] vreg_48_3;
	node n48_3(.left(vreg_47_3), .right(vreg_49_3), .up(vreg_48_4), .down(vreg_48_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_3), .sw(sw));
	wire signed[17:0] vwire_48_4;
	reg signed[17:0] vreg_48_4;
	node n48_4(.left(vreg_47_4), .right(vreg_49_4), .up(vreg_48_5), .down(vreg_48_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_4), .sw(sw));
	wire signed[17:0] vwire_48_5;
	reg signed[17:0] vreg_48_5;
	node n48_5(.left(vreg_47_5), .right(vreg_49_5), .up(vreg_48_6), .down(vreg_48_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_5), .sw(sw));
	wire signed[17:0] vwire_48_6;
	reg signed[17:0] vreg_48_6;
	node n48_6(.left(vreg_47_6), .right(vreg_49_6), .up(vreg_48_7), .down(vreg_48_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_6), .sw(sw));
	wire signed[17:0] vwire_48_7;
	reg signed[17:0] vreg_48_7;
	node n48_7(.left(vreg_47_7), .right(vreg_49_7), .up(vreg_48_8), .down(vreg_48_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_7), .sw(sw));
	wire signed[17:0] vwire_48_8;
	reg signed[17:0] vreg_48_8;
	node n48_8(.left(vreg_47_8), .right(vreg_49_8), .up(vreg_48_9), .down(vreg_48_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_8), .sw(sw));
	wire signed[17:0] vwire_48_9;
	reg signed[17:0] vreg_48_9;
	node n48_9(.left(vreg_47_9), .right(vreg_49_9), .up(vreg_48_10), .down(vreg_48_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_9), .sw(sw));
	wire signed[17:0] vwire_48_10;
	reg signed[17:0] vreg_48_10;
	node n48_10(.left(vreg_47_10), .right(vreg_49_10), .up(vreg_48_11), .down(vreg_48_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_10), .sw(sw));
	wire signed[17:0] vwire_48_11;
	reg signed[17:0] vreg_48_11;
	node n48_11(.left(vreg_47_11), .right(vreg_49_11), .up(vreg_48_12), .down(vreg_48_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_11), .sw(sw));
	wire signed[17:0] vwire_48_12;
	reg signed[17:0] vreg_48_12;
	node n48_12(.left(vreg_47_12), .right(vreg_49_12), .up(vreg_48_13), .down(vreg_48_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_12), .sw(sw));
	wire signed[17:0] vwire_48_13;
	reg signed[17:0] vreg_48_13;
	node n48_13(.left(vreg_47_13), .right(vreg_49_13), .up(vreg_48_14), .down(vreg_48_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_13), .sw(sw));
	wire signed[17:0] vwire_48_14;
	reg signed[17:0] vreg_48_14;
	node n48_14(.left(vreg_47_14), .right(vreg_49_14), .up(vreg_48_15), .down(vreg_48_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_14), .sw(sw));
	wire signed[17:0] vwire_48_15;
	reg signed[17:0] vreg_48_15;
	node n48_15(.left(vreg_47_15), .right(vreg_49_15), .up(vreg_48_16), .down(vreg_48_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_15), .sw(sw));
	wire signed[17:0] vwire_48_16;
	reg signed[17:0] vreg_48_16;
	node n48_16(.left(vreg_47_16), .right(vreg_49_16), .up(vreg_48_17), .down(vreg_48_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_16), .sw(sw));
	wire signed[17:0] vwire_48_17;
	reg signed[17:0] vreg_48_17;
	node n48_17(.left(vreg_47_17), .right(vreg_49_17), .up(vreg_48_18), .down(vreg_48_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_17), .sw(sw));
	wire signed[17:0] vwire_48_18;
	reg signed[17:0] vreg_48_18;
	node n48_18(.left(vreg_47_18), .right(vreg_49_18), .up(vreg_48_19), .down(vreg_48_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_18), .sw(sw));
	wire signed[17:0] vwire_48_19;
	reg signed[17:0] vreg_48_19;
	node n48_19(.left(vreg_47_19), .right(vreg_49_19), .up(vreg_48_20), .down(vreg_48_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_19), .sw(sw));
	wire signed[17:0] vwire_48_20;
	reg signed[17:0] vreg_48_20;
	node n48_20(.left(vreg_47_20), .right(vreg_49_20), .up(vreg_48_21), .down(vreg_48_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_20), .sw(sw));
	wire signed[17:0] vwire_48_21;
	reg signed[17:0] vreg_48_21;
	node n48_21(.left(vreg_47_21), .right(vreg_49_21), .up(vreg_48_22), .down(vreg_48_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_21), .sw(sw));
	wire signed[17:0] vwire_48_22;
	reg signed[17:0] vreg_48_22;
	node n48_22(.left(vreg_47_22), .right(vreg_49_22), .up(vreg_48_23), .down(vreg_48_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_22), .sw(sw));
	wire signed[17:0] vwire_48_23;
	reg signed[17:0] vreg_48_23;
	node n48_23(.left(vreg_47_23), .right(vreg_49_23), .up(vreg_48_24), .down(vreg_48_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_23), .sw(sw));
	wire signed[17:0] vwire_48_24;
	reg signed[17:0] vreg_48_24;
	node n48_24(.left(vreg_47_24), .right(vreg_49_24), .up(vreg_48_25), .down(vreg_48_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_24), .sw(sw));
	wire signed[17:0] vwire_48_25;
	reg signed[17:0] vreg_48_25;
	node n48_25(.left(vreg_47_25), .right(vreg_49_25), .up(vreg_48_26), .down(vreg_48_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_25), .sw(sw));
	wire signed[17:0] vwire_48_26;
	reg signed[17:0] vreg_48_26;
	node n48_26(.left(vreg_47_26), .right(vreg_49_26), .up(vreg_48_27), .down(vreg_48_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_26), .sw(sw));
	wire signed[17:0] vwire_48_27;
	reg signed[17:0] vreg_48_27;
	node n48_27(.left(vreg_47_27), .right(vreg_49_27), .up(vreg_48_28), .down(vreg_48_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_27), .sw(sw));
	wire signed[17:0] vwire_48_28;
	reg signed[17:0] vreg_48_28;
	node n48_28(.left(vreg_47_28), .right(vreg_49_28), .up(vreg_48_29), .down(vreg_48_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_28), .sw(sw));
	wire signed[17:0] vwire_48_29;
	reg signed[17:0] vreg_48_29;
	node n48_29(.left(vreg_47_29), .right(vreg_49_29), .up(vreg_48_30), .down(vreg_48_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_29), .sw(sw));
	wire signed[17:0] vwire_48_30;
	reg signed[17:0] vreg_48_30;
	node n48_30(.left(vreg_47_30), .right(vreg_49_30), .up(vreg_48_31), .down(vreg_48_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_30), .sw(sw));
	wire signed[17:0] vwire_48_31;
	reg signed[17:0] vreg_48_31;
	node n48_31(.left(vreg_47_31), .right(vreg_49_31), .up(vreg_48_32), .down(vreg_48_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_31), .sw(sw));
	wire signed[17:0] vwire_48_32;
	reg signed[17:0] vreg_48_32;
	node n48_32(.left(vreg_47_32), .right(vreg_49_32), .up(vreg_48_33), .down(vreg_48_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_32), .sw(sw));
	wire signed[17:0] vwire_48_33;
	reg signed[17:0] vreg_48_33;
	node n48_33(.left(vreg_47_33), .right(vreg_49_33), .up(vreg_48_34), .down(vreg_48_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_33), .sw(sw));
	wire signed[17:0] vwire_48_34;
	reg signed[17:0] vreg_48_34;
	node n48_34(.left(vreg_47_34), .right(vreg_49_34), .up(vreg_48_35), .down(vreg_48_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_34), .sw(sw));
	wire signed[17:0] vwire_48_35;
	reg signed[17:0] vreg_48_35;
	node n48_35(.left(vreg_47_35), .right(vreg_49_35), .up(vreg_48_36), .down(vreg_48_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_35), .sw(sw));
	wire signed[17:0] vwire_48_36;
	reg signed[17:0] vreg_48_36;
	node n48_36(.left(vreg_47_36), .right(vreg_49_36), .up(vreg_48_37), .down(vreg_48_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_36), .sw(sw));
	wire signed[17:0] vwire_48_37;
	reg signed[17:0] vreg_48_37;
	node n48_37(.left(vreg_47_37), .right(vreg_49_37), .up(vreg_48_38), .down(vreg_48_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_37), .sw(sw));
	wire signed[17:0] vwire_48_38;
	reg signed[17:0] vreg_48_38;
	node n48_38(.left(vreg_47_38), .right(vreg_49_38), .up(vreg_48_39), .down(vreg_48_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_38), .sw(sw));
	wire signed[17:0] vwire_48_39;
	reg signed[17:0] vreg_48_39;
	node n48_39(.left(vreg_47_39), .right(vreg_49_39), .up(vreg_48_40), .down(vreg_48_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_39), .sw(sw));
	wire signed[17:0] vwire_48_40;
	reg signed[17:0] vreg_48_40;
	node n48_40(.left(vreg_47_40), .right(vreg_49_40), .up(vreg_48_41), .down(vreg_48_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_40), .sw(sw));
	wire signed[17:0] vwire_48_41;
	reg signed[17:0] vreg_48_41;
	node n48_41(.left(vreg_47_41), .right(vreg_49_41), .up(vreg_48_42), .down(vreg_48_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_41), .sw(sw));
	wire signed[17:0] vwire_48_42;
	reg signed[17:0] vreg_48_42;
	node n48_42(.left(vreg_47_42), .right(vreg_49_42), .up(vreg_48_43), .down(vreg_48_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_42), .sw(sw));
	wire signed[17:0] vwire_48_43;
	reg signed[17:0] vreg_48_43;
	node n48_43(.left(vreg_47_43), .right(vreg_49_43), .up(vreg_48_44), .down(vreg_48_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_43), .sw(sw));
	wire signed[17:0] vwire_48_44;
	reg signed[17:0] vreg_48_44;
	node n48_44(.left(vreg_47_44), .right(vreg_49_44), .up(vreg_48_45), .down(vreg_48_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_44), .sw(sw));
	wire signed[17:0] vwire_48_45;
	reg signed[17:0] vreg_48_45;
	node n48_45(.left(vreg_47_45), .right(vreg_49_45), .up(vreg_48_46), .down(vreg_48_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_45), .sw(sw));
	wire signed[17:0] vwire_48_46;
	reg signed[17:0] vreg_48_46;
	node n48_46(.left(vreg_47_46), .right(vreg_49_46), .up(vreg_48_47), .down(vreg_48_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_46), .sw(sw));
	wire signed[17:0] vwire_48_47;
	reg signed[17:0] vreg_48_47;
	node n48_47(.left(vreg_47_47), .right(vreg_49_47), .up(vreg_48_48), .down(vreg_48_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_47), .sw(sw));
	wire signed[17:0] vwire_48_48;
	reg signed[17:0] vreg_48_48;
	node n48_48(.left(vreg_47_48), .right(vreg_49_48), .up(vreg_48_49), .down(vreg_48_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_48), .sw(sw));
	wire signed[17:0] vwire_48_49;
	reg signed[17:0] vreg_48_49;
	node n48_49(.left(vreg_47_49), .right(vreg_49_49), .up(18'b0), .down(vreg_48_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_48_49), .sw(sw));
	wire signed[17:0] vwire_49_0;
	reg signed[17:0] vreg_49_0;
	node n49_0(.left(vreg_48_0), .right(18'b0), .up(vreg_49_1), .down(vreg_49_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_0), .sw(sw));
	wire signed[17:0] vwire_49_1;
	reg signed[17:0] vreg_49_1;
	node n49_1(.left(vreg_48_1), .right(18'b0), .up(vreg_49_2), .down(vreg_49_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_1), .sw(sw));
	wire signed[17:0] vwire_49_2;
	reg signed[17:0] vreg_49_2;
	node n49_2(.left(vreg_48_2), .right(18'b0), .up(vreg_49_3), .down(vreg_49_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_2), .sw(sw));
	wire signed[17:0] vwire_49_3;
	reg signed[17:0] vreg_49_3;
	node n49_3(.left(vreg_48_3), .right(18'b0), .up(vreg_49_4), .down(vreg_49_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_3), .sw(sw));
	wire signed[17:0] vwire_49_4;
	reg signed[17:0] vreg_49_4;
	node n49_4(.left(vreg_48_4), .right(18'b0), .up(vreg_49_5), .down(vreg_49_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_4), .sw(sw));
	wire signed[17:0] vwire_49_5;
	reg signed[17:0] vreg_49_5;
	node n49_5(.left(vreg_48_5), .right(18'b0), .up(vreg_49_6), .down(vreg_49_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_5), .sw(sw));
	wire signed[17:0] vwire_49_6;
	reg signed[17:0] vreg_49_6;
	node n49_6(.left(vreg_48_6), .right(18'b0), .up(vreg_49_7), .down(vreg_49_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_6), .sw(sw));
	wire signed[17:0] vwire_49_7;
	reg signed[17:0] vreg_49_7;
	node n49_7(.left(vreg_48_7), .right(18'b0), .up(vreg_49_8), .down(vreg_49_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_7), .sw(sw));
	wire signed[17:0] vwire_49_8;
	reg signed[17:0] vreg_49_8;
	node n49_8(.left(vreg_48_8), .right(18'b0), .up(vreg_49_9), .down(vreg_49_7), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_8), .sw(sw));
	wire signed[17:0] vwire_49_9;
	reg signed[17:0] vreg_49_9;
	node n49_9(.left(vreg_48_9), .right(18'b0), .up(vreg_49_10), .down(vreg_49_8), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_9), .sw(sw));
	wire signed[17:0] vwire_49_10;
	reg signed[17:0] vreg_49_10;
	node n49_10(.left(vreg_48_10), .right(18'b0), .up(vreg_49_11), .down(vreg_49_9), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_10), .sw(sw));
	wire signed[17:0] vwire_49_11;
	reg signed[17:0] vreg_49_11;
	node n49_11(.left(vreg_48_11), .right(18'b0), .up(vreg_49_12), .down(vreg_49_10), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_11), .sw(sw));
	wire signed[17:0] vwire_49_12;
	reg signed[17:0] vreg_49_12;
	node n49_12(.left(vreg_48_12), .right(18'b0), .up(vreg_49_13), .down(vreg_49_11), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_12), .sw(sw));
	wire signed[17:0] vwire_49_13;
	reg signed[17:0] vreg_49_13;
	node n49_13(.left(vreg_48_13), .right(18'b0), .up(vreg_49_14), .down(vreg_49_12), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_13), .sw(sw));
	wire signed[17:0] vwire_49_14;
	reg signed[17:0] vreg_49_14;
	node n49_14(.left(vreg_48_14), .right(18'b0), .up(vreg_49_15), .down(vreg_49_13), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_14), .sw(sw));
	wire signed[17:0] vwire_49_15;
	reg signed[17:0] vreg_49_15;
	node n49_15(.left(vreg_48_15), .right(18'b0), .up(vreg_49_16), .down(vreg_49_14), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_15), .sw(sw));
	wire signed[17:0] vwire_49_16;
	reg signed[17:0] vreg_49_16;
	node n49_16(.left(vreg_48_16), .right(18'b0), .up(vreg_49_17), .down(vreg_49_15), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_16), .sw(sw));
	wire signed[17:0] vwire_49_17;
	reg signed[17:0] vreg_49_17;
	node n49_17(.left(vreg_48_17), .right(18'b0), .up(vreg_49_18), .down(vreg_49_16), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_17), .sw(sw));
	wire signed[17:0] vwire_49_18;
	reg signed[17:0] vreg_49_18;
	node n49_18(.left(vreg_48_18), .right(18'b0), .up(vreg_49_19), .down(vreg_49_17), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_18), .sw(sw));
	wire signed[17:0] vwire_49_19;
	reg signed[17:0] vreg_49_19;
	node n49_19(.left(vreg_48_19), .right(18'b0), .up(vreg_49_20), .down(vreg_49_18), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_19), .sw(sw));
	wire signed[17:0] vwire_49_20;
	reg signed[17:0] vreg_49_20;
	node n49_20(.left(vreg_48_20), .right(18'b0), .up(vreg_49_21), .down(vreg_49_19), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_20), .sw(sw));
	wire signed[17:0] vwire_49_21;
	reg signed[17:0] vreg_49_21;
	node n49_21(.left(vreg_48_21), .right(18'b0), .up(vreg_49_22), .down(vreg_49_20), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_21), .sw(sw));
	wire signed[17:0] vwire_49_22;
	reg signed[17:0] vreg_49_22;
	node n49_22(.left(vreg_48_22), .right(18'b0), .up(vreg_49_23), .down(vreg_49_21), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_22), .sw(sw));
	wire signed[17:0] vwire_49_23;
	reg signed[17:0] vreg_49_23;
	node n49_23(.left(vreg_48_23), .right(18'b0), .up(vreg_49_24), .down(vreg_49_22), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_23), .sw(sw));
	wire signed[17:0] vwire_49_24;
	reg signed[17:0] vreg_49_24;
	node n49_24(.left(vreg_48_24), .right(18'b0), .up(vreg_49_25), .down(vreg_49_23), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_24), .sw(sw));
	wire signed[17:0] vwire_49_25;
	reg signed[17:0] vreg_49_25;
	node n49_25(.left(vreg_48_25), .right(18'b0), .up(vreg_49_26), .down(vreg_49_24), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_25), .sw(sw));
	wire signed[17:0] vwire_49_26;
	reg signed[17:0] vreg_49_26;
	node n49_26(.left(vreg_48_26), .right(18'b0), .up(vreg_49_27), .down(vreg_49_25), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_26), .sw(sw));
	wire signed[17:0] vwire_49_27;
	reg signed[17:0] vreg_49_27;
	node n49_27(.left(vreg_48_27), .right(18'b0), .up(vreg_49_28), .down(vreg_49_26), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_27), .sw(sw));
	wire signed[17:0] vwire_49_28;
	reg signed[17:0] vreg_49_28;
	node n49_28(.left(vreg_48_28), .right(18'b0), .up(vreg_49_29), .down(vreg_49_27), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_28), .sw(sw));
	wire signed[17:0] vwire_49_29;
	reg signed[17:0] vreg_49_29;
	node n49_29(.left(vreg_48_29), .right(18'b0), .up(vreg_49_30), .down(vreg_49_28), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_29), .sw(sw));
	wire signed[17:0] vwire_49_30;
	reg signed[17:0] vreg_49_30;
	node n49_30(.left(vreg_48_30), .right(18'b0), .up(vreg_49_31), .down(vreg_49_29), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_30), .sw(sw));
	wire signed[17:0] vwire_49_31;
	reg signed[17:0] vreg_49_31;
	node n49_31(.left(vreg_48_31), .right(18'b0), .up(vreg_49_32), .down(vreg_49_30), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_31), .sw(sw));
	wire signed[17:0] vwire_49_32;
	reg signed[17:0] vreg_49_32;
	node n49_32(.left(vreg_48_32), .right(18'b0), .up(vreg_49_33), .down(vreg_49_31), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_32), .sw(sw));
	wire signed[17:0] vwire_49_33;
	reg signed[17:0] vreg_49_33;
	node n49_33(.left(vreg_48_33), .right(18'b0), .up(vreg_49_34), .down(vreg_49_32), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_33), .sw(sw));
	wire signed[17:0] vwire_49_34;
	reg signed[17:0] vreg_49_34;
	node n49_34(.left(vreg_48_34), .right(18'b0), .up(vreg_49_35), .down(vreg_49_33), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_34), .sw(sw));
	wire signed[17:0] vwire_49_35;
	reg signed[17:0] vreg_49_35;
	node n49_35(.left(vreg_48_35), .right(18'b0), .up(vreg_49_36), .down(vreg_49_34), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_35), .sw(sw));
	wire signed[17:0] vwire_49_36;
	reg signed[17:0] vreg_49_36;
	node n49_36(.left(vreg_48_36), .right(18'b0), .up(vreg_49_37), .down(vreg_49_35), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_36), .sw(sw));
	wire signed[17:0] vwire_49_37;
	reg signed[17:0] vreg_49_37;
	node n49_37(.left(vreg_48_37), .right(18'b0), .up(vreg_49_38), .down(vreg_49_36), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_37), .sw(sw));
	wire signed[17:0] vwire_49_38;
	reg signed[17:0] vreg_49_38;
	node n49_38(.left(vreg_48_38), .right(18'b0), .up(vreg_49_39), .down(vreg_49_37), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_38), .sw(sw));
	wire signed[17:0] vwire_49_39;
	reg signed[17:0] vreg_49_39;
	node n49_39(.left(vreg_48_39), .right(18'b0), .up(vreg_49_40), .down(vreg_49_38), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_39), .sw(sw));
	wire signed[17:0] vwire_49_40;
	reg signed[17:0] vreg_49_40;
	node n49_40(.left(vreg_48_40), .right(18'b0), .up(vreg_49_41), .down(vreg_49_39), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_40), .sw(sw));
	wire signed[17:0] vwire_49_41;
	reg signed[17:0] vreg_49_41;
	node n49_41(.left(vreg_48_41), .right(18'b0), .up(vreg_49_42), .down(vreg_49_40), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_41), .sw(sw));
	wire signed[17:0] vwire_49_42;
	reg signed[17:0] vreg_49_42;
	node n49_42(.left(vreg_48_42), .right(18'b0), .up(vreg_49_43), .down(vreg_49_41), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_42), .sw(sw));
	wire signed[17:0] vwire_49_43;
	reg signed[17:0] vreg_49_43;
	node n49_43(.left(vreg_48_43), .right(18'b0), .up(vreg_49_44), .down(vreg_49_42), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_43), .sw(sw));
	wire signed[17:0] vwire_49_44;
	reg signed[17:0] vreg_49_44;
	node n49_44(.left(vreg_48_44), .right(18'b0), .up(vreg_49_45), .down(vreg_49_43), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_44), .sw(sw));
	wire signed[17:0] vwire_49_45;
	reg signed[17:0] vreg_49_45;
	node n49_45(.left(vreg_48_45), .right(18'b0), .up(vreg_49_46), .down(vreg_49_44), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_45), .sw(sw));
	wire signed[17:0] vwire_49_46;
	reg signed[17:0] vreg_49_46;
	node n49_46(.left(vreg_48_46), .right(18'b0), .up(vreg_49_47), .down(vreg_49_45), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_46), .sw(sw));
	wire signed[17:0] vwire_49_47;
	reg signed[17:0] vreg_49_47;
	node n49_47(.left(vreg_48_47), .right(18'b0), .up(vreg_49_48), .down(vreg_49_46), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_47), .sw(sw));
	wire signed[17:0] vwire_49_48;
	reg signed[17:0] vreg_49_48;
	node n49_48(.left(vreg_48_48), .right(18'b0), .up(vreg_49_49), .down(vreg_49_47), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_48), .sw(sw));
	wire signed[17:0] vwire_49_49;
	reg signed[17:0] vreg_49_49;
	node n49_49(.left(vreg_48_49), .right(18'b0), .up(18'b0), .down(vreg_49_48), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_49_49), .sw(sw));
	always @ (negedge clk)
	begin
		vreg_0_0 <= vwire_0_0;
		vreg_0_1 <= vwire_0_1;
		vreg_0_2 <= vwire_0_2;
		vreg_0_3 <= vwire_0_3;
		vreg_0_4 <= vwire_0_4;
		vreg_0_5 <= vwire_0_5;
		vreg_0_6 <= vwire_0_6;
		vreg_0_7 <= vwire_0_7;
		vreg_0_8 <= vwire_0_8;
		vreg_0_9 <= vwire_0_9;
		vreg_0_10 <= vwire_0_10;
		vreg_0_11 <= vwire_0_11;
		vreg_0_12 <= vwire_0_12;
		vreg_0_13 <= vwire_0_13;
		vreg_0_14 <= vwire_0_14;
		vreg_0_15 <= vwire_0_15;
		vreg_0_16 <= vwire_0_16;
		vreg_0_17 <= vwire_0_17;
		vreg_0_18 <= vwire_0_18;
		vreg_0_19 <= vwire_0_19;
		vreg_0_20 <= vwire_0_20;
		vreg_0_21 <= vwire_0_21;
		vreg_0_22 <= vwire_0_22;
		vreg_0_23 <= vwire_0_23;
		vreg_0_24 <= vwire_0_24;
		vreg_0_25 <= vwire_0_25;
		vreg_0_26 <= vwire_0_26;
		vreg_0_27 <= vwire_0_27;
		vreg_0_28 <= vwire_0_28;
		vreg_0_29 <= vwire_0_29;
		vreg_0_30 <= vwire_0_30;
		vreg_0_31 <= vwire_0_31;
		vreg_0_32 <= vwire_0_32;
		vreg_0_33 <= vwire_0_33;
		vreg_0_34 <= vwire_0_34;
		vreg_0_35 <= vwire_0_35;
		vreg_0_36 <= vwire_0_36;
		vreg_0_37 <= vwire_0_37;
		vreg_0_38 <= vwire_0_38;
		vreg_0_39 <= vwire_0_39;
		vreg_0_40 <= vwire_0_40;
		vreg_0_41 <= vwire_0_41;
		vreg_0_42 <= vwire_0_42;
		vreg_0_43 <= vwire_0_43;
		vreg_0_44 <= vwire_0_44;
		vreg_0_45 <= vwire_0_45;
		vreg_0_46 <= vwire_0_46;
		vreg_0_47 <= vwire_0_47;
		vreg_0_48 <= vwire_0_48;
		vreg_0_49 <= vwire_0_49;
		vreg_1_0 <= vwire_1_0;
		vreg_1_1 <= vwire_1_1;
		vreg_1_2 <= vwire_1_2;
		vreg_1_3 <= vwire_1_3;
		vreg_1_4 <= vwire_1_4;
		vreg_1_5 <= vwire_1_5;
		vreg_1_6 <= vwire_1_6;
		vreg_1_7 <= vwire_1_7;
		vreg_1_8 <= vwire_1_8;
		vreg_1_9 <= vwire_1_9;
		vreg_1_10 <= vwire_1_10;
		vreg_1_11 <= vwire_1_11;
		vreg_1_12 <= vwire_1_12;
		vreg_1_13 <= vwire_1_13;
		vreg_1_14 <= vwire_1_14;
		vreg_1_15 <= vwire_1_15;
		vreg_1_16 <= vwire_1_16;
		vreg_1_17 <= vwire_1_17;
		vreg_1_18 <= vwire_1_18;
		vreg_1_19 <= vwire_1_19;
		vreg_1_20 <= vwire_1_20;
		vreg_1_21 <= vwire_1_21;
		vreg_1_22 <= vwire_1_22;
		vreg_1_23 <= vwire_1_23;
		vreg_1_24 <= vwire_1_24;
		vreg_1_25 <= vwire_1_25;
		vreg_1_26 <= vwire_1_26;
		vreg_1_27 <= vwire_1_27;
		vreg_1_28 <= vwire_1_28;
		vreg_1_29 <= vwire_1_29;
		vreg_1_30 <= vwire_1_30;
		vreg_1_31 <= vwire_1_31;
		vreg_1_32 <= vwire_1_32;
		vreg_1_33 <= vwire_1_33;
		vreg_1_34 <= vwire_1_34;
		vreg_1_35 <= vwire_1_35;
		vreg_1_36 <= vwire_1_36;
		vreg_1_37 <= vwire_1_37;
		vreg_1_38 <= vwire_1_38;
		vreg_1_39 <= vwire_1_39;
		vreg_1_40 <= vwire_1_40;
		vreg_1_41 <= vwire_1_41;
		vreg_1_42 <= vwire_1_42;
		vreg_1_43 <= vwire_1_43;
		vreg_1_44 <= vwire_1_44;
		vreg_1_45 <= vwire_1_45;
		vreg_1_46 <= vwire_1_46;
		vreg_1_47 <= vwire_1_47;
		vreg_1_48 <= vwire_1_48;
		vreg_1_49 <= vwire_1_49;
		vreg_2_0 <= vwire_2_0;
		vreg_2_1 <= vwire_2_1;
		vreg_2_2 <= vwire_2_2;
		vreg_2_3 <= vwire_2_3;
		vreg_2_4 <= vwire_2_4;
		vreg_2_5 <= vwire_2_5;
		vreg_2_6 <= vwire_2_6;
		vreg_2_7 <= vwire_2_7;
		vreg_2_8 <= vwire_2_8;
		vreg_2_9 <= vwire_2_9;
		vreg_2_10 <= vwire_2_10;
		vreg_2_11 <= vwire_2_11;
		vreg_2_12 <= vwire_2_12;
		vreg_2_13 <= vwire_2_13;
		vreg_2_14 <= vwire_2_14;
		vreg_2_15 <= vwire_2_15;
		vreg_2_16 <= vwire_2_16;
		vreg_2_17 <= vwire_2_17;
		vreg_2_18 <= vwire_2_18;
		vreg_2_19 <= vwire_2_19;
		vreg_2_20 <= vwire_2_20;
		vreg_2_21 <= vwire_2_21;
		vreg_2_22 <= vwire_2_22;
		vreg_2_23 <= vwire_2_23;
		vreg_2_24 <= vwire_2_24;
		vreg_2_25 <= vwire_2_25;
		vreg_2_26 <= vwire_2_26;
		vreg_2_27 <= vwire_2_27;
		vreg_2_28 <= vwire_2_28;
		vreg_2_29 <= vwire_2_29;
		vreg_2_30 <= vwire_2_30;
		vreg_2_31 <= vwire_2_31;
		vreg_2_32 <= vwire_2_32;
		vreg_2_33 <= vwire_2_33;
		vreg_2_34 <= vwire_2_34;
		vreg_2_35 <= vwire_2_35;
		vreg_2_36 <= vwire_2_36;
		vreg_2_37 <= vwire_2_37;
		vreg_2_38 <= vwire_2_38;
		vreg_2_39 <= vwire_2_39;
		vreg_2_40 <= vwire_2_40;
		vreg_2_41 <= vwire_2_41;
		vreg_2_42 <= vwire_2_42;
		vreg_2_43 <= vwire_2_43;
		vreg_2_44 <= vwire_2_44;
		vreg_2_45 <= vwire_2_45;
		vreg_2_46 <= vwire_2_46;
		vreg_2_47 <= vwire_2_47;
		vreg_2_48 <= vwire_2_48;
		vreg_2_49 <= vwire_2_49;
		vreg_3_0 <= vwire_3_0;
		vreg_3_1 <= vwire_3_1;
		vreg_3_2 <= vwire_3_2;
		vreg_3_3 <= vwire_3_3;
		vreg_3_4 <= vwire_3_4;
		vreg_3_5 <= vwire_3_5;
		vreg_3_6 <= vwire_3_6;
		vreg_3_7 <= vwire_3_7;
		vreg_3_8 <= vwire_3_8;
		vreg_3_9 <= vwire_3_9;
		vreg_3_10 <= vwire_3_10;
		vreg_3_11 <= vwire_3_11;
		vreg_3_12 <= vwire_3_12;
		vreg_3_13 <= vwire_3_13;
		vreg_3_14 <= vwire_3_14;
		vreg_3_15 <= vwire_3_15;
		vreg_3_16 <= vwire_3_16;
		vreg_3_17 <= vwire_3_17;
		vreg_3_18 <= vwire_3_18;
		vreg_3_19 <= vwire_3_19;
		vreg_3_20 <= vwire_3_20;
		vreg_3_21 <= vwire_3_21;
		vreg_3_22 <= vwire_3_22;
		vreg_3_23 <= vwire_3_23;
		vreg_3_24 <= vwire_3_24;
		vreg_3_25 <= vwire_3_25;
		vreg_3_26 <= vwire_3_26;
		vreg_3_27 <= vwire_3_27;
		vreg_3_28 <= vwire_3_28;
		vreg_3_29 <= vwire_3_29;
		vreg_3_30 <= vwire_3_30;
		vreg_3_31 <= vwire_3_31;
		vreg_3_32 <= vwire_3_32;
		vreg_3_33 <= vwire_3_33;
		vreg_3_34 <= vwire_3_34;
		vreg_3_35 <= vwire_3_35;
		vreg_3_36 <= vwire_3_36;
		vreg_3_37 <= vwire_3_37;
		vreg_3_38 <= vwire_3_38;
		vreg_3_39 <= vwire_3_39;
		vreg_3_40 <= vwire_3_40;
		vreg_3_41 <= vwire_3_41;
		vreg_3_42 <= vwire_3_42;
		vreg_3_43 <= vwire_3_43;
		vreg_3_44 <= vwire_3_44;
		vreg_3_45 <= vwire_3_45;
		vreg_3_46 <= vwire_3_46;
		vreg_3_47 <= vwire_3_47;
		vreg_3_48 <= vwire_3_48;
		vreg_3_49 <= vwire_3_49;
		vreg_4_0 <= vwire_4_0;
		vreg_4_1 <= vwire_4_1;
		vreg_4_2 <= vwire_4_2;
		vreg_4_3 <= vwire_4_3;
		vreg_4_4 <= vwire_4_4;
		vreg_4_5 <= vwire_4_5;
		vreg_4_6 <= vwire_4_6;
		vreg_4_7 <= vwire_4_7;
		vreg_4_8 <= vwire_4_8;
		vreg_4_9 <= vwire_4_9;
		vreg_4_10 <= vwire_4_10;
		vreg_4_11 <= vwire_4_11;
		vreg_4_12 <= vwire_4_12;
		vreg_4_13 <= vwire_4_13;
		vreg_4_14 <= vwire_4_14;
		vreg_4_15 <= vwire_4_15;
		vreg_4_16 <= vwire_4_16;
		vreg_4_17 <= vwire_4_17;
		vreg_4_18 <= vwire_4_18;
		vreg_4_19 <= vwire_4_19;
		vreg_4_20 <= vwire_4_20;
		vreg_4_21 <= vwire_4_21;
		vreg_4_22 <= vwire_4_22;
		vreg_4_23 <= vwire_4_23;
		vreg_4_24 <= vwire_4_24;
		vreg_4_25 <= vwire_4_25;
		vreg_4_26 <= vwire_4_26;
		vreg_4_27 <= vwire_4_27;
		vreg_4_28 <= vwire_4_28;
		vreg_4_29 <= vwire_4_29;
		vreg_4_30 <= vwire_4_30;
		vreg_4_31 <= vwire_4_31;
		vreg_4_32 <= vwire_4_32;
		vreg_4_33 <= vwire_4_33;
		vreg_4_34 <= vwire_4_34;
		vreg_4_35 <= vwire_4_35;
		vreg_4_36 <= vwire_4_36;
		vreg_4_37 <= vwire_4_37;
		vreg_4_38 <= vwire_4_38;
		vreg_4_39 <= vwire_4_39;
		vreg_4_40 <= vwire_4_40;
		vreg_4_41 <= vwire_4_41;
		vreg_4_42 <= vwire_4_42;
		vreg_4_43 <= vwire_4_43;
		vreg_4_44 <= vwire_4_44;
		vreg_4_45 <= vwire_4_45;
		vreg_4_46 <= vwire_4_46;
		vreg_4_47 <= vwire_4_47;
		vreg_4_48 <= vwire_4_48;
		vreg_4_49 <= vwire_4_49;
		vreg_5_0 <= vwire_5_0;
		vreg_5_1 <= vwire_5_1;
		vreg_5_2 <= vwire_5_2;
		vreg_5_3 <= vwire_5_3;
		vreg_5_4 <= vwire_5_4;
		vreg_5_5 <= vwire_5_5;
		vreg_5_6 <= vwire_5_6;
		vreg_5_7 <= vwire_5_7;
		vreg_5_8 <= vwire_5_8;
		vreg_5_9 <= vwire_5_9;
		vreg_5_10 <= vwire_5_10;
		vreg_5_11 <= vwire_5_11;
		vreg_5_12 <= vwire_5_12;
		vreg_5_13 <= vwire_5_13;
		vreg_5_14 <= vwire_5_14;
		vreg_5_15 <= vwire_5_15;
		vreg_5_16 <= vwire_5_16;
		vreg_5_17 <= vwire_5_17;
		vreg_5_18 <= vwire_5_18;
		vreg_5_19 <= vwire_5_19;
		vreg_5_20 <= vwire_5_20;
		vreg_5_21 <= vwire_5_21;
		vreg_5_22 <= vwire_5_22;
		vreg_5_23 <= vwire_5_23;
		vreg_5_24 <= vwire_5_24;
		vreg_5_25 <= vwire_5_25;
		vreg_5_26 <= vwire_5_26;
		vreg_5_27 <= vwire_5_27;
		vreg_5_28 <= vwire_5_28;
		vreg_5_29 <= vwire_5_29;
		vreg_5_30 <= vwire_5_30;
		vreg_5_31 <= vwire_5_31;
		vreg_5_32 <= vwire_5_32;
		vreg_5_33 <= vwire_5_33;
		vreg_5_34 <= vwire_5_34;
		vreg_5_35 <= vwire_5_35;
		vreg_5_36 <= vwire_5_36;
		vreg_5_37 <= vwire_5_37;
		vreg_5_38 <= vwire_5_38;
		vreg_5_39 <= vwire_5_39;
		vreg_5_40 <= vwire_5_40;
		vreg_5_41 <= vwire_5_41;
		vreg_5_42 <= vwire_5_42;
		vreg_5_43 <= vwire_5_43;
		vreg_5_44 <= vwire_5_44;
		vreg_5_45 <= vwire_5_45;
		vreg_5_46 <= vwire_5_46;
		vreg_5_47 <= vwire_5_47;
		vreg_5_48 <= vwire_5_48;
		vreg_5_49 <= vwire_5_49;
		vreg_6_0 <= vwire_6_0;
		vreg_6_1 <= vwire_6_1;
		vreg_6_2 <= vwire_6_2;
		vreg_6_3 <= vwire_6_3;
		vreg_6_4 <= vwire_6_4;
		vreg_6_5 <= vwire_6_5;
		vreg_6_6 <= vwire_6_6;
		vreg_6_7 <= vwire_6_7;
		vreg_6_8 <= vwire_6_8;
		vreg_6_9 <= vwire_6_9;
		vreg_6_10 <= vwire_6_10;
		vreg_6_11 <= vwire_6_11;
		vreg_6_12 <= vwire_6_12;
		vreg_6_13 <= vwire_6_13;
		vreg_6_14 <= vwire_6_14;
		vreg_6_15 <= vwire_6_15;
		vreg_6_16 <= vwire_6_16;
		vreg_6_17 <= vwire_6_17;
		vreg_6_18 <= vwire_6_18;
		vreg_6_19 <= vwire_6_19;
		vreg_6_20 <= vwire_6_20;
		vreg_6_21 <= vwire_6_21;
		vreg_6_22 <= vwire_6_22;
		vreg_6_23 <= vwire_6_23;
		vreg_6_24 <= vwire_6_24;
		vreg_6_25 <= vwire_6_25;
		vreg_6_26 <= vwire_6_26;
		vreg_6_27 <= vwire_6_27;
		vreg_6_28 <= vwire_6_28;
		vreg_6_29 <= vwire_6_29;
		vreg_6_30 <= vwire_6_30;
		vreg_6_31 <= vwire_6_31;
		vreg_6_32 <= vwire_6_32;
		vreg_6_33 <= vwire_6_33;
		vreg_6_34 <= vwire_6_34;
		vreg_6_35 <= vwire_6_35;
		vreg_6_36 <= vwire_6_36;
		vreg_6_37 <= vwire_6_37;
		vreg_6_38 <= vwire_6_38;
		vreg_6_39 <= vwire_6_39;
		vreg_6_40 <= vwire_6_40;
		vreg_6_41 <= vwire_6_41;
		vreg_6_42 <= vwire_6_42;
		vreg_6_43 <= vwire_6_43;
		vreg_6_44 <= vwire_6_44;
		vreg_6_45 <= vwire_6_45;
		vreg_6_46 <= vwire_6_46;
		vreg_6_47 <= vwire_6_47;
		vreg_6_48 <= vwire_6_48;
		vreg_6_49 <= vwire_6_49;
		vreg_7_0 <= vwire_7_0;
		vreg_7_1 <= vwire_7_1;
		vreg_7_2 <= vwire_7_2;
		vreg_7_3 <= vwire_7_3;
		vreg_7_4 <= vwire_7_4;
		vreg_7_5 <= vwire_7_5;
		vreg_7_6 <= vwire_7_6;
		vreg_7_7 <= vwire_7_7;
		vreg_7_8 <= vwire_7_8;
		vreg_7_9 <= vwire_7_9;
		vreg_7_10 <= vwire_7_10;
		vreg_7_11 <= vwire_7_11;
		vreg_7_12 <= vwire_7_12;
		vreg_7_13 <= vwire_7_13;
		vreg_7_14 <= vwire_7_14;
		vreg_7_15 <= vwire_7_15;
		vreg_7_16 <= vwire_7_16;
		vreg_7_17 <= vwire_7_17;
		vreg_7_18 <= vwire_7_18;
		vreg_7_19 <= vwire_7_19;
		vreg_7_20 <= vwire_7_20;
		vreg_7_21 <= vwire_7_21;
		vreg_7_22 <= vwire_7_22;
		vreg_7_23 <= vwire_7_23;
		vreg_7_24 <= vwire_7_24;
		vreg_7_25 <= vwire_7_25;
		vreg_7_26 <= vwire_7_26;
		vreg_7_27 <= vwire_7_27;
		vreg_7_28 <= vwire_7_28;
		vreg_7_29 <= vwire_7_29;
		vreg_7_30 <= vwire_7_30;
		vreg_7_31 <= vwire_7_31;
		vreg_7_32 <= vwire_7_32;
		vreg_7_33 <= vwire_7_33;
		vreg_7_34 <= vwire_7_34;
		vreg_7_35 <= vwire_7_35;
		vreg_7_36 <= vwire_7_36;
		vreg_7_37 <= vwire_7_37;
		vreg_7_38 <= vwire_7_38;
		vreg_7_39 <= vwire_7_39;
		vreg_7_40 <= vwire_7_40;
		vreg_7_41 <= vwire_7_41;
		vreg_7_42 <= vwire_7_42;
		vreg_7_43 <= vwire_7_43;
		vreg_7_44 <= vwire_7_44;
		vreg_7_45 <= vwire_7_45;
		vreg_7_46 <= vwire_7_46;
		vreg_7_47 <= vwire_7_47;
		vreg_7_48 <= vwire_7_48;
		vreg_7_49 <= vwire_7_49;
		vreg_8_0 <= vwire_8_0;
		vreg_8_1 <= vwire_8_1;
		vreg_8_2 <= vwire_8_2;
		vreg_8_3 <= vwire_8_3;
		vreg_8_4 <= vwire_8_4;
		vreg_8_5 <= vwire_8_5;
		vreg_8_6 <= vwire_8_6;
		vreg_8_7 <= vwire_8_7;
		vreg_8_8 <= vwire_8_8;
		vreg_8_9 <= vwire_8_9;
		vreg_8_10 <= vwire_8_10;
		vreg_8_11 <= vwire_8_11;
		vreg_8_12 <= vwire_8_12;
		vreg_8_13 <= vwire_8_13;
		vreg_8_14 <= vwire_8_14;
		vreg_8_15 <= vwire_8_15;
		vreg_8_16 <= vwire_8_16;
		vreg_8_17 <= vwire_8_17;
		vreg_8_18 <= vwire_8_18;
		vreg_8_19 <= vwire_8_19;
		vreg_8_20 <= vwire_8_20;
		vreg_8_21 <= vwire_8_21;
		vreg_8_22 <= vwire_8_22;
		vreg_8_23 <= vwire_8_23;
		vreg_8_24 <= vwire_8_24;
		vreg_8_25 <= vwire_8_25;
		vreg_8_26 <= vwire_8_26;
		vreg_8_27 <= vwire_8_27;
		vreg_8_28 <= vwire_8_28;
		vreg_8_29 <= vwire_8_29;
		vreg_8_30 <= vwire_8_30;
		vreg_8_31 <= vwire_8_31;
		vreg_8_32 <= vwire_8_32;
		vreg_8_33 <= vwire_8_33;
		vreg_8_34 <= vwire_8_34;
		vreg_8_35 <= vwire_8_35;
		vreg_8_36 <= vwire_8_36;
		vreg_8_37 <= vwire_8_37;
		vreg_8_38 <= vwire_8_38;
		vreg_8_39 <= vwire_8_39;
		vreg_8_40 <= vwire_8_40;
		vreg_8_41 <= vwire_8_41;
		vreg_8_42 <= vwire_8_42;
		vreg_8_43 <= vwire_8_43;
		vreg_8_44 <= vwire_8_44;
		vreg_8_45 <= vwire_8_45;
		vreg_8_46 <= vwire_8_46;
		vreg_8_47 <= vwire_8_47;
		vreg_8_48 <= vwire_8_48;
		vreg_8_49 <= vwire_8_49;
		vreg_9_0 <= vwire_9_0;
		vreg_9_1 <= vwire_9_1;
		vreg_9_2 <= vwire_9_2;
		vreg_9_3 <= vwire_9_3;
		vreg_9_4 <= vwire_9_4;
		vreg_9_5 <= vwire_9_5;
		vreg_9_6 <= vwire_9_6;
		vreg_9_7 <= vwire_9_7;
		vreg_9_8 <= vwire_9_8;
		vreg_9_9 <= vwire_9_9;
		vreg_9_10 <= vwire_9_10;
		vreg_9_11 <= vwire_9_11;
		vreg_9_12 <= vwire_9_12;
		vreg_9_13 <= vwire_9_13;
		vreg_9_14 <= vwire_9_14;
		vreg_9_15 <= vwire_9_15;
		vreg_9_16 <= vwire_9_16;
		vreg_9_17 <= vwire_9_17;
		vreg_9_18 <= vwire_9_18;
		vreg_9_19 <= vwire_9_19;
		vreg_9_20 <= vwire_9_20;
		vreg_9_21 <= vwire_9_21;
		vreg_9_22 <= vwire_9_22;
		vreg_9_23 <= vwire_9_23;
		vreg_9_24 <= vwire_9_24;
		vreg_9_25 <= vwire_9_25;
		vreg_9_26 <= vwire_9_26;
		vreg_9_27 <= vwire_9_27;
		vreg_9_28 <= vwire_9_28;
		vreg_9_29 <= vwire_9_29;
		vreg_9_30 <= vwire_9_30;
		vreg_9_31 <= vwire_9_31;
		vreg_9_32 <= vwire_9_32;
		vreg_9_33 <= vwire_9_33;
		vreg_9_34 <= vwire_9_34;
		vreg_9_35 <= vwire_9_35;
		vreg_9_36 <= vwire_9_36;
		vreg_9_37 <= vwire_9_37;
		vreg_9_38 <= vwire_9_38;
		vreg_9_39 <= vwire_9_39;
		vreg_9_40 <= vwire_9_40;
		vreg_9_41 <= vwire_9_41;
		vreg_9_42 <= vwire_9_42;
		vreg_9_43 <= vwire_9_43;
		vreg_9_44 <= vwire_9_44;
		vreg_9_45 <= vwire_9_45;
		vreg_9_46 <= vwire_9_46;
		vreg_9_47 <= vwire_9_47;
		vreg_9_48 <= vwire_9_48;
		vreg_9_49 <= vwire_9_49;
		vreg_10_0 <= vwire_10_0;
		vreg_10_1 <= vwire_10_1;
		vreg_10_2 <= vwire_10_2;
		vreg_10_3 <= vwire_10_3;
		vreg_10_4 <= vwire_10_4;
		vreg_10_5 <= vwire_10_5;
		vreg_10_6 <= vwire_10_6;
		vreg_10_7 <= vwire_10_7;
		vreg_10_8 <= vwire_10_8;
		vreg_10_9 <= vwire_10_9;
		vreg_10_10 <= vwire_10_10;
		vreg_10_11 <= vwire_10_11;
		vreg_10_12 <= vwire_10_12;
		vreg_10_13 <= vwire_10_13;
		vreg_10_14 <= vwire_10_14;
		vreg_10_15 <= vwire_10_15;
		vreg_10_16 <= vwire_10_16;
		vreg_10_17 <= vwire_10_17;
		vreg_10_18 <= vwire_10_18;
		vreg_10_19 <= vwire_10_19;
		vreg_10_20 <= vwire_10_20;
		vreg_10_21 <= vwire_10_21;
		vreg_10_22 <= vwire_10_22;
		vreg_10_23 <= vwire_10_23;
		vreg_10_24 <= vwire_10_24;
		vreg_10_25 <= vwire_10_25;
		vreg_10_26 <= vwire_10_26;
		vreg_10_27 <= vwire_10_27;
		vreg_10_28 <= vwire_10_28;
		vreg_10_29 <= vwire_10_29;
		vreg_10_30 <= vwire_10_30;
		vreg_10_31 <= vwire_10_31;
		vreg_10_32 <= vwire_10_32;
		vreg_10_33 <= vwire_10_33;
		vreg_10_34 <= vwire_10_34;
		vreg_10_35 <= vwire_10_35;
		vreg_10_36 <= vwire_10_36;
		vreg_10_37 <= vwire_10_37;
		vreg_10_38 <= vwire_10_38;
		vreg_10_39 <= vwire_10_39;
		vreg_10_40 <= vwire_10_40;
		vreg_10_41 <= vwire_10_41;
		vreg_10_42 <= vwire_10_42;
		vreg_10_43 <= vwire_10_43;
		vreg_10_44 <= vwire_10_44;
		vreg_10_45 <= vwire_10_45;
		vreg_10_46 <= vwire_10_46;
		vreg_10_47 <= vwire_10_47;
		vreg_10_48 <= vwire_10_48;
		vreg_10_49 <= vwire_10_49;
		vreg_11_0 <= vwire_11_0;
		vreg_11_1 <= vwire_11_1;
		vreg_11_2 <= vwire_11_2;
		vreg_11_3 <= vwire_11_3;
		vreg_11_4 <= vwire_11_4;
		vreg_11_5 <= vwire_11_5;
		vreg_11_6 <= vwire_11_6;
		vreg_11_7 <= vwire_11_7;
		vreg_11_8 <= vwire_11_8;
		vreg_11_9 <= vwire_11_9;
		vreg_11_10 <= vwire_11_10;
		vreg_11_11 <= vwire_11_11;
		vreg_11_12 <= vwire_11_12;
		vreg_11_13 <= vwire_11_13;
		vreg_11_14 <= vwire_11_14;
		vreg_11_15 <= vwire_11_15;
		vreg_11_16 <= vwire_11_16;
		vreg_11_17 <= vwire_11_17;
		vreg_11_18 <= vwire_11_18;
		vreg_11_19 <= vwire_11_19;
		vreg_11_20 <= vwire_11_20;
		vreg_11_21 <= vwire_11_21;
		vreg_11_22 <= vwire_11_22;
		vreg_11_23 <= vwire_11_23;
		vreg_11_24 <= vwire_11_24;
		vreg_11_25 <= vwire_11_25;
		vreg_11_26 <= vwire_11_26;
		vreg_11_27 <= vwire_11_27;
		vreg_11_28 <= vwire_11_28;
		vreg_11_29 <= vwire_11_29;
		vreg_11_30 <= vwire_11_30;
		vreg_11_31 <= vwire_11_31;
		vreg_11_32 <= vwire_11_32;
		vreg_11_33 <= vwire_11_33;
		vreg_11_34 <= vwire_11_34;
		vreg_11_35 <= vwire_11_35;
		vreg_11_36 <= vwire_11_36;
		vreg_11_37 <= vwire_11_37;
		vreg_11_38 <= vwire_11_38;
		vreg_11_39 <= vwire_11_39;
		vreg_11_40 <= vwire_11_40;
		vreg_11_41 <= vwire_11_41;
		vreg_11_42 <= vwire_11_42;
		vreg_11_43 <= vwire_11_43;
		vreg_11_44 <= vwire_11_44;
		vreg_11_45 <= vwire_11_45;
		vreg_11_46 <= vwire_11_46;
		vreg_11_47 <= vwire_11_47;
		vreg_11_48 <= vwire_11_48;
		vreg_11_49 <= vwire_11_49;
		vreg_12_0 <= vwire_12_0;
		vreg_12_1 <= vwire_12_1;
		vreg_12_2 <= vwire_12_2;
		vreg_12_3 <= vwire_12_3;
		vreg_12_4 <= vwire_12_4;
		vreg_12_5 <= vwire_12_5;
		vreg_12_6 <= vwire_12_6;
		vreg_12_7 <= vwire_12_7;
		vreg_12_8 <= vwire_12_8;
		vreg_12_9 <= vwire_12_9;
		vreg_12_10 <= vwire_12_10;
		vreg_12_11 <= vwire_12_11;
		vreg_12_12 <= vwire_12_12;
		vreg_12_13 <= vwire_12_13;
		vreg_12_14 <= vwire_12_14;
		vreg_12_15 <= vwire_12_15;
		vreg_12_16 <= vwire_12_16;
		vreg_12_17 <= vwire_12_17;
		vreg_12_18 <= vwire_12_18;
		vreg_12_19 <= vwire_12_19;
		vreg_12_20 <= vwire_12_20;
		vreg_12_21 <= vwire_12_21;
		vreg_12_22 <= vwire_12_22;
		vreg_12_23 <= vwire_12_23;
		vreg_12_24 <= vwire_12_24;
		vreg_12_25 <= vwire_12_25;
		vreg_12_26 <= vwire_12_26;
		vreg_12_27 <= vwire_12_27;
		vreg_12_28 <= vwire_12_28;
		vreg_12_29 <= vwire_12_29;
		vreg_12_30 <= vwire_12_30;
		vreg_12_31 <= vwire_12_31;
		vreg_12_32 <= vwire_12_32;
		vreg_12_33 <= vwire_12_33;
		vreg_12_34 <= vwire_12_34;
		vreg_12_35 <= vwire_12_35;
		vreg_12_36 <= vwire_12_36;
		vreg_12_37 <= vwire_12_37;
		vreg_12_38 <= vwire_12_38;
		vreg_12_39 <= vwire_12_39;
		vreg_12_40 <= vwire_12_40;
		vreg_12_41 <= vwire_12_41;
		vreg_12_42 <= vwire_12_42;
		vreg_12_43 <= vwire_12_43;
		vreg_12_44 <= vwire_12_44;
		vreg_12_45 <= vwire_12_45;
		vreg_12_46 <= vwire_12_46;
		vreg_12_47 <= vwire_12_47;
		vreg_12_48 <= vwire_12_48;
		vreg_12_49 <= vwire_12_49;
		vreg_13_0 <= vwire_13_0;
		vreg_13_1 <= vwire_13_1;
		vreg_13_2 <= vwire_13_2;
		vreg_13_3 <= vwire_13_3;
		vreg_13_4 <= vwire_13_4;
		vreg_13_5 <= vwire_13_5;
		vreg_13_6 <= vwire_13_6;
		vreg_13_7 <= vwire_13_7;
		vreg_13_8 <= vwire_13_8;
		vreg_13_9 <= vwire_13_9;
		vreg_13_10 <= vwire_13_10;
		vreg_13_11 <= vwire_13_11;
		vreg_13_12 <= vwire_13_12;
		vreg_13_13 <= vwire_13_13;
		vreg_13_14 <= vwire_13_14;
		vreg_13_15 <= vwire_13_15;
		vreg_13_16 <= vwire_13_16;
		vreg_13_17 <= vwire_13_17;
		vreg_13_18 <= vwire_13_18;
		vreg_13_19 <= vwire_13_19;
		vreg_13_20 <= vwire_13_20;
		vreg_13_21 <= vwire_13_21;
		vreg_13_22 <= vwire_13_22;
		vreg_13_23 <= vwire_13_23;
		vreg_13_24 <= vwire_13_24;
		vreg_13_25 <= vwire_13_25;
		vreg_13_26 <= vwire_13_26;
		vreg_13_27 <= vwire_13_27;
		vreg_13_28 <= vwire_13_28;
		vreg_13_29 <= vwire_13_29;
		vreg_13_30 <= vwire_13_30;
		vreg_13_31 <= vwire_13_31;
		vreg_13_32 <= vwire_13_32;
		vreg_13_33 <= vwire_13_33;
		vreg_13_34 <= vwire_13_34;
		vreg_13_35 <= vwire_13_35;
		vreg_13_36 <= vwire_13_36;
		vreg_13_37 <= vwire_13_37;
		vreg_13_38 <= vwire_13_38;
		vreg_13_39 <= vwire_13_39;
		vreg_13_40 <= vwire_13_40;
		vreg_13_41 <= vwire_13_41;
		vreg_13_42 <= vwire_13_42;
		vreg_13_43 <= vwire_13_43;
		vreg_13_44 <= vwire_13_44;
		vreg_13_45 <= vwire_13_45;
		vreg_13_46 <= vwire_13_46;
		vreg_13_47 <= vwire_13_47;
		vreg_13_48 <= vwire_13_48;
		vreg_13_49 <= vwire_13_49;
		vreg_14_0 <= vwire_14_0;
		vreg_14_1 <= vwire_14_1;
		vreg_14_2 <= vwire_14_2;
		vreg_14_3 <= vwire_14_3;
		vreg_14_4 <= vwire_14_4;
		vreg_14_5 <= vwire_14_5;
		vreg_14_6 <= vwire_14_6;
		vreg_14_7 <= vwire_14_7;
		vreg_14_8 <= vwire_14_8;
		vreg_14_9 <= vwire_14_9;
		vreg_14_10 <= vwire_14_10;
		vreg_14_11 <= vwire_14_11;
		vreg_14_12 <= vwire_14_12;
		vreg_14_13 <= vwire_14_13;
		vreg_14_14 <= vwire_14_14;
		vreg_14_15 <= vwire_14_15;
		vreg_14_16 <= vwire_14_16;
		vreg_14_17 <= vwire_14_17;
		vreg_14_18 <= vwire_14_18;
		vreg_14_19 <= vwire_14_19;
		vreg_14_20 <= vwire_14_20;
		vreg_14_21 <= vwire_14_21;
		vreg_14_22 <= vwire_14_22;
		vreg_14_23 <= vwire_14_23;
		vreg_14_24 <= vwire_14_24;
		vreg_14_25 <= vwire_14_25;
		vreg_14_26 <= vwire_14_26;
		vreg_14_27 <= vwire_14_27;
		vreg_14_28 <= vwire_14_28;
		vreg_14_29 <= vwire_14_29;
		vreg_14_30 <= vwire_14_30;
		vreg_14_31 <= vwire_14_31;
		vreg_14_32 <= vwire_14_32;
		vreg_14_33 <= vwire_14_33;
		vreg_14_34 <= vwire_14_34;
		vreg_14_35 <= vwire_14_35;
		vreg_14_36 <= vwire_14_36;
		vreg_14_37 <= vwire_14_37;
		vreg_14_38 <= vwire_14_38;
		vreg_14_39 <= vwire_14_39;
		vreg_14_40 <= vwire_14_40;
		vreg_14_41 <= vwire_14_41;
		vreg_14_42 <= vwire_14_42;
		vreg_14_43 <= vwire_14_43;
		vreg_14_44 <= vwire_14_44;
		vreg_14_45 <= vwire_14_45;
		vreg_14_46 <= vwire_14_46;
		vreg_14_47 <= vwire_14_47;
		vreg_14_48 <= vwire_14_48;
		vreg_14_49 <= vwire_14_49;
		vreg_15_0 <= vwire_15_0;
		vreg_15_1 <= vwire_15_1;
		vreg_15_2 <= vwire_15_2;
		vreg_15_3 <= vwire_15_3;
		vreg_15_4 <= vwire_15_4;
		vreg_15_5 <= vwire_15_5;
		vreg_15_6 <= vwire_15_6;
		vreg_15_7 <= vwire_15_7;
		vreg_15_8 <= vwire_15_8;
		vreg_15_9 <= vwire_15_9;
		vreg_15_10 <= vwire_15_10;
		vreg_15_11 <= vwire_15_11;
		vreg_15_12 <= vwire_15_12;
		vreg_15_13 <= vwire_15_13;
		vreg_15_14 <= vwire_15_14;
		vreg_15_15 <= vwire_15_15;
		vreg_15_16 <= vwire_15_16;
		vreg_15_17 <= vwire_15_17;
		vreg_15_18 <= vwire_15_18;
		vreg_15_19 <= vwire_15_19;
		vreg_15_20 <= vwire_15_20;
		vreg_15_21 <= vwire_15_21;
		vreg_15_22 <= vwire_15_22;
		vreg_15_23 <= vwire_15_23;
		vreg_15_24 <= vwire_15_24;
		vreg_15_25 <= vwire_15_25;
		vreg_15_26 <= vwire_15_26;
		vreg_15_27 <= vwire_15_27;
		vreg_15_28 <= vwire_15_28;
		vreg_15_29 <= vwire_15_29;
		vreg_15_30 <= vwire_15_30;
		vreg_15_31 <= vwire_15_31;
		vreg_15_32 <= vwire_15_32;
		vreg_15_33 <= vwire_15_33;
		vreg_15_34 <= vwire_15_34;
		vreg_15_35 <= vwire_15_35;
		vreg_15_36 <= vwire_15_36;
		vreg_15_37 <= vwire_15_37;
		vreg_15_38 <= vwire_15_38;
		vreg_15_39 <= vwire_15_39;
		vreg_15_40 <= vwire_15_40;
		vreg_15_41 <= vwire_15_41;
		vreg_15_42 <= vwire_15_42;
		vreg_15_43 <= vwire_15_43;
		vreg_15_44 <= vwire_15_44;
		vreg_15_45 <= vwire_15_45;
		vreg_15_46 <= vwire_15_46;
		vreg_15_47 <= vwire_15_47;
		vreg_15_48 <= vwire_15_48;
		vreg_15_49 <= vwire_15_49;
		vreg_16_0 <= vwire_16_0;
		vreg_16_1 <= vwire_16_1;
		vreg_16_2 <= vwire_16_2;
		vreg_16_3 <= vwire_16_3;
		vreg_16_4 <= vwire_16_4;
		vreg_16_5 <= vwire_16_5;
		vreg_16_6 <= vwire_16_6;
		vreg_16_7 <= vwire_16_7;
		vreg_16_8 <= vwire_16_8;
		vreg_16_9 <= vwire_16_9;
		vreg_16_10 <= vwire_16_10;
		vreg_16_11 <= vwire_16_11;
		vreg_16_12 <= vwire_16_12;
		vreg_16_13 <= vwire_16_13;
		vreg_16_14 <= vwire_16_14;
		vreg_16_15 <= vwire_16_15;
		vreg_16_16 <= vwire_16_16;
		vreg_16_17 <= vwire_16_17;
		vreg_16_18 <= vwire_16_18;
		vreg_16_19 <= vwire_16_19;
		vreg_16_20 <= vwire_16_20;
		vreg_16_21 <= vwire_16_21;
		vreg_16_22 <= vwire_16_22;
		vreg_16_23 <= vwire_16_23;
		vreg_16_24 <= vwire_16_24;
		vreg_16_25 <= vwire_16_25;
		vreg_16_26 <= vwire_16_26;
		vreg_16_27 <= vwire_16_27;
		vreg_16_28 <= vwire_16_28;
		vreg_16_29 <= vwire_16_29;
		vreg_16_30 <= vwire_16_30;
		vreg_16_31 <= vwire_16_31;
		vreg_16_32 <= vwire_16_32;
		vreg_16_33 <= vwire_16_33;
		vreg_16_34 <= vwire_16_34;
		vreg_16_35 <= vwire_16_35;
		vreg_16_36 <= vwire_16_36;
		vreg_16_37 <= vwire_16_37;
		vreg_16_38 <= vwire_16_38;
		vreg_16_39 <= vwire_16_39;
		vreg_16_40 <= vwire_16_40;
		vreg_16_41 <= vwire_16_41;
		vreg_16_42 <= vwire_16_42;
		vreg_16_43 <= vwire_16_43;
		vreg_16_44 <= vwire_16_44;
		vreg_16_45 <= vwire_16_45;
		vreg_16_46 <= vwire_16_46;
		vreg_16_47 <= vwire_16_47;
		vreg_16_48 <= vwire_16_48;
		vreg_16_49 <= vwire_16_49;
		vreg_17_0 <= vwire_17_0;
		vreg_17_1 <= vwire_17_1;
		vreg_17_2 <= vwire_17_2;
		vreg_17_3 <= vwire_17_3;
		vreg_17_4 <= vwire_17_4;
		vreg_17_5 <= vwire_17_5;
		vreg_17_6 <= vwire_17_6;
		vreg_17_7 <= vwire_17_7;
		vreg_17_8 <= vwire_17_8;
		vreg_17_9 <= vwire_17_9;
		vreg_17_10 <= vwire_17_10;
		vreg_17_11 <= vwire_17_11;
		vreg_17_12 <= vwire_17_12;
		vreg_17_13 <= vwire_17_13;
		vreg_17_14 <= vwire_17_14;
		vreg_17_15 <= vwire_17_15;
		vreg_17_16 <= vwire_17_16;
		vreg_17_17 <= vwire_17_17;
		vreg_17_18 <= vwire_17_18;
		vreg_17_19 <= vwire_17_19;
		vreg_17_20 <= vwire_17_20;
		vreg_17_21 <= vwire_17_21;
		vreg_17_22 <= vwire_17_22;
		vreg_17_23 <= vwire_17_23;
		vreg_17_24 <= vwire_17_24;
		vreg_17_25 <= vwire_17_25;
		vreg_17_26 <= vwire_17_26;
		vreg_17_27 <= vwire_17_27;
		vreg_17_28 <= vwire_17_28;
		vreg_17_29 <= vwire_17_29;
		vreg_17_30 <= vwire_17_30;
		vreg_17_31 <= vwire_17_31;
		vreg_17_32 <= vwire_17_32;
		vreg_17_33 <= vwire_17_33;
		vreg_17_34 <= vwire_17_34;
		vreg_17_35 <= vwire_17_35;
		vreg_17_36 <= vwire_17_36;
		vreg_17_37 <= vwire_17_37;
		vreg_17_38 <= vwire_17_38;
		vreg_17_39 <= vwire_17_39;
		vreg_17_40 <= vwire_17_40;
		vreg_17_41 <= vwire_17_41;
		vreg_17_42 <= vwire_17_42;
		vreg_17_43 <= vwire_17_43;
		vreg_17_44 <= vwire_17_44;
		vreg_17_45 <= vwire_17_45;
		vreg_17_46 <= vwire_17_46;
		vreg_17_47 <= vwire_17_47;
		vreg_17_48 <= vwire_17_48;
		vreg_17_49 <= vwire_17_49;
		vreg_18_0 <= vwire_18_0;
		vreg_18_1 <= vwire_18_1;
		vreg_18_2 <= vwire_18_2;
		vreg_18_3 <= vwire_18_3;
		vreg_18_4 <= vwire_18_4;
		vreg_18_5 <= vwire_18_5;
		vreg_18_6 <= vwire_18_6;
		vreg_18_7 <= vwire_18_7;
		vreg_18_8 <= vwire_18_8;
		vreg_18_9 <= vwire_18_9;
		vreg_18_10 <= vwire_18_10;
		vreg_18_11 <= vwire_18_11;
		vreg_18_12 <= vwire_18_12;
		vreg_18_13 <= vwire_18_13;
		vreg_18_14 <= vwire_18_14;
		vreg_18_15 <= vwire_18_15;
		vreg_18_16 <= vwire_18_16;
		vreg_18_17 <= vwire_18_17;
		vreg_18_18 <= vwire_18_18;
		vreg_18_19 <= vwire_18_19;
		vreg_18_20 <= vwire_18_20;
		vreg_18_21 <= vwire_18_21;
		vreg_18_22 <= vwire_18_22;
		vreg_18_23 <= vwire_18_23;
		vreg_18_24 <= vwire_18_24;
		vreg_18_25 <= vwire_18_25;
		vreg_18_26 <= vwire_18_26;
		vreg_18_27 <= vwire_18_27;
		vreg_18_28 <= vwire_18_28;
		vreg_18_29 <= vwire_18_29;
		vreg_18_30 <= vwire_18_30;
		vreg_18_31 <= vwire_18_31;
		vreg_18_32 <= vwire_18_32;
		vreg_18_33 <= vwire_18_33;
		vreg_18_34 <= vwire_18_34;
		vreg_18_35 <= vwire_18_35;
		vreg_18_36 <= vwire_18_36;
		vreg_18_37 <= vwire_18_37;
		vreg_18_38 <= vwire_18_38;
		vreg_18_39 <= vwire_18_39;
		vreg_18_40 <= vwire_18_40;
		vreg_18_41 <= vwire_18_41;
		vreg_18_42 <= vwire_18_42;
		vreg_18_43 <= vwire_18_43;
		vreg_18_44 <= vwire_18_44;
		vreg_18_45 <= vwire_18_45;
		vreg_18_46 <= vwire_18_46;
		vreg_18_47 <= vwire_18_47;
		vreg_18_48 <= vwire_18_48;
		vreg_18_49 <= vwire_18_49;
		vreg_19_0 <= vwire_19_0;
		vreg_19_1 <= vwire_19_1;
		vreg_19_2 <= vwire_19_2;
		vreg_19_3 <= vwire_19_3;
		vreg_19_4 <= vwire_19_4;
		vreg_19_5 <= vwire_19_5;
		vreg_19_6 <= vwire_19_6;
		vreg_19_7 <= vwire_19_7;
		vreg_19_8 <= vwire_19_8;
		vreg_19_9 <= vwire_19_9;
		vreg_19_10 <= vwire_19_10;
		vreg_19_11 <= vwire_19_11;
		vreg_19_12 <= vwire_19_12;
		vreg_19_13 <= vwire_19_13;
		vreg_19_14 <= vwire_19_14;
		vreg_19_15 <= vwire_19_15;
		vreg_19_16 <= vwire_19_16;
		vreg_19_17 <= vwire_19_17;
		vreg_19_18 <= vwire_19_18;
		vreg_19_19 <= vwire_19_19;
		vreg_19_20 <= vwire_19_20;
		vreg_19_21 <= vwire_19_21;
		vreg_19_22 <= vwire_19_22;
		vreg_19_23 <= vwire_19_23;
		vreg_19_24 <= vwire_19_24;
		vreg_19_25 <= vwire_19_25;
		vreg_19_26 <= vwire_19_26;
		vreg_19_27 <= vwire_19_27;
		vreg_19_28 <= vwire_19_28;
		vreg_19_29 <= vwire_19_29;
		vreg_19_30 <= vwire_19_30;
		vreg_19_31 <= vwire_19_31;
		vreg_19_32 <= vwire_19_32;
		vreg_19_33 <= vwire_19_33;
		vreg_19_34 <= vwire_19_34;
		vreg_19_35 <= vwire_19_35;
		vreg_19_36 <= vwire_19_36;
		vreg_19_37 <= vwire_19_37;
		vreg_19_38 <= vwire_19_38;
		vreg_19_39 <= vwire_19_39;
		vreg_19_40 <= vwire_19_40;
		vreg_19_41 <= vwire_19_41;
		vreg_19_42 <= vwire_19_42;
		vreg_19_43 <= vwire_19_43;
		vreg_19_44 <= vwire_19_44;
		vreg_19_45 <= vwire_19_45;
		vreg_19_46 <= vwire_19_46;
		vreg_19_47 <= vwire_19_47;
		vreg_19_48 <= vwire_19_48;
		vreg_19_49 <= vwire_19_49;
		vreg_20_0 <= vwire_20_0;
		vreg_20_1 <= vwire_20_1;
		vreg_20_2 <= vwire_20_2;
		vreg_20_3 <= vwire_20_3;
		vreg_20_4 <= vwire_20_4;
		vreg_20_5 <= vwire_20_5;
		vreg_20_6 <= vwire_20_6;
		vreg_20_7 <= vwire_20_7;
		vreg_20_8 <= vwire_20_8;
		vreg_20_9 <= vwire_20_9;
		vreg_20_10 <= vwire_20_10;
		vreg_20_11 <= vwire_20_11;
		vreg_20_12 <= vwire_20_12;
		vreg_20_13 <= vwire_20_13;
		vreg_20_14 <= vwire_20_14;
		vreg_20_15 <= vwire_20_15;
		vreg_20_16 <= vwire_20_16;
		vreg_20_17 <= vwire_20_17;
		vreg_20_18 <= vwire_20_18;
		vreg_20_19 <= vwire_20_19;
		vreg_20_20 <= vwire_20_20;
		vreg_20_21 <= vwire_20_21;
		vreg_20_22 <= vwire_20_22;
		vreg_20_23 <= vwire_20_23;
		vreg_20_24 <= vwire_20_24;
		vreg_20_25 <= vwire_20_25;
		vreg_20_26 <= vwire_20_26;
		vreg_20_27 <= vwire_20_27;
		vreg_20_28 <= vwire_20_28;
		vreg_20_29 <= vwire_20_29;
		vreg_20_30 <= vwire_20_30;
		vreg_20_31 <= vwire_20_31;
		vreg_20_32 <= vwire_20_32;
		vreg_20_33 <= vwire_20_33;
		vreg_20_34 <= vwire_20_34;
		vreg_20_35 <= vwire_20_35;
		vreg_20_36 <= vwire_20_36;
		vreg_20_37 <= vwire_20_37;
		vreg_20_38 <= vwire_20_38;
		vreg_20_39 <= vwire_20_39;
		vreg_20_40 <= vwire_20_40;
		vreg_20_41 <= vwire_20_41;
		vreg_20_42 <= vwire_20_42;
		vreg_20_43 <= vwire_20_43;
		vreg_20_44 <= vwire_20_44;
		vreg_20_45 <= vwire_20_45;
		vreg_20_46 <= vwire_20_46;
		vreg_20_47 <= vwire_20_47;
		vreg_20_48 <= vwire_20_48;
		vreg_20_49 <= vwire_20_49;
		vreg_21_0 <= vwire_21_0;
		vreg_21_1 <= vwire_21_1;
		vreg_21_2 <= vwire_21_2;
		vreg_21_3 <= vwire_21_3;
		vreg_21_4 <= vwire_21_4;
		vreg_21_5 <= vwire_21_5;
		vreg_21_6 <= vwire_21_6;
		vreg_21_7 <= vwire_21_7;
		vreg_21_8 <= vwire_21_8;
		vreg_21_9 <= vwire_21_9;
		vreg_21_10 <= vwire_21_10;
		vreg_21_11 <= vwire_21_11;
		vreg_21_12 <= vwire_21_12;
		vreg_21_13 <= vwire_21_13;
		vreg_21_14 <= vwire_21_14;
		vreg_21_15 <= vwire_21_15;
		vreg_21_16 <= vwire_21_16;
		vreg_21_17 <= vwire_21_17;
		vreg_21_18 <= vwire_21_18;
		vreg_21_19 <= vwire_21_19;
		vreg_21_20 <= vwire_21_20;
		vreg_21_21 <= vwire_21_21;
		vreg_21_22 <= vwire_21_22;
		vreg_21_23 <= vwire_21_23;
		vreg_21_24 <= vwire_21_24;
		vreg_21_25 <= vwire_21_25;
		vreg_21_26 <= vwire_21_26;
		vreg_21_27 <= vwire_21_27;
		vreg_21_28 <= vwire_21_28;
		vreg_21_29 <= vwire_21_29;
		vreg_21_30 <= vwire_21_30;
		vreg_21_31 <= vwire_21_31;
		vreg_21_32 <= vwire_21_32;
		vreg_21_33 <= vwire_21_33;
		vreg_21_34 <= vwire_21_34;
		vreg_21_35 <= vwire_21_35;
		vreg_21_36 <= vwire_21_36;
		vreg_21_37 <= vwire_21_37;
		vreg_21_38 <= vwire_21_38;
		vreg_21_39 <= vwire_21_39;
		vreg_21_40 <= vwire_21_40;
		vreg_21_41 <= vwire_21_41;
		vreg_21_42 <= vwire_21_42;
		vreg_21_43 <= vwire_21_43;
		vreg_21_44 <= vwire_21_44;
		vreg_21_45 <= vwire_21_45;
		vreg_21_46 <= vwire_21_46;
		vreg_21_47 <= vwire_21_47;
		vreg_21_48 <= vwire_21_48;
		vreg_21_49 <= vwire_21_49;
		vreg_22_0 <= vwire_22_0;
		vreg_22_1 <= vwire_22_1;
		vreg_22_2 <= vwire_22_2;
		vreg_22_3 <= vwire_22_3;
		vreg_22_4 <= vwire_22_4;
		vreg_22_5 <= vwire_22_5;
		vreg_22_6 <= vwire_22_6;
		vreg_22_7 <= vwire_22_7;
		vreg_22_8 <= vwire_22_8;
		vreg_22_9 <= vwire_22_9;
		vreg_22_10 <= vwire_22_10;
		vreg_22_11 <= vwire_22_11;
		vreg_22_12 <= vwire_22_12;
		vreg_22_13 <= vwire_22_13;
		vreg_22_14 <= vwire_22_14;
		vreg_22_15 <= vwire_22_15;
		vreg_22_16 <= vwire_22_16;
		vreg_22_17 <= vwire_22_17;
		vreg_22_18 <= vwire_22_18;
		vreg_22_19 <= vwire_22_19;
		vreg_22_20 <= vwire_22_20;
		vreg_22_21 <= vwire_22_21;
		vreg_22_22 <= vwire_22_22;
		vreg_22_23 <= vwire_22_23;
		vreg_22_24 <= vwire_22_24;
		vreg_22_25 <= vwire_22_25;
		vreg_22_26 <= vwire_22_26;
		vreg_22_27 <= vwire_22_27;
		vreg_22_28 <= vwire_22_28;
		vreg_22_29 <= vwire_22_29;
		vreg_22_30 <= vwire_22_30;
		vreg_22_31 <= vwire_22_31;
		vreg_22_32 <= vwire_22_32;
		vreg_22_33 <= vwire_22_33;
		vreg_22_34 <= vwire_22_34;
		vreg_22_35 <= vwire_22_35;
		vreg_22_36 <= vwire_22_36;
		vreg_22_37 <= vwire_22_37;
		vreg_22_38 <= vwire_22_38;
		vreg_22_39 <= vwire_22_39;
		vreg_22_40 <= vwire_22_40;
		vreg_22_41 <= vwire_22_41;
		vreg_22_42 <= vwire_22_42;
		vreg_22_43 <= vwire_22_43;
		vreg_22_44 <= vwire_22_44;
		vreg_22_45 <= vwire_22_45;
		vreg_22_46 <= vwire_22_46;
		vreg_22_47 <= vwire_22_47;
		vreg_22_48 <= vwire_22_48;
		vreg_22_49 <= vwire_22_49;
		vreg_23_0 <= vwire_23_0;
		vreg_23_1 <= vwire_23_1;
		vreg_23_2 <= vwire_23_2;
		vreg_23_3 <= vwire_23_3;
		vreg_23_4 <= vwire_23_4;
		vreg_23_5 <= vwire_23_5;
		vreg_23_6 <= vwire_23_6;
		vreg_23_7 <= vwire_23_7;
		vreg_23_8 <= vwire_23_8;
		vreg_23_9 <= vwire_23_9;
		vreg_23_10 <= vwire_23_10;
		vreg_23_11 <= vwire_23_11;
		vreg_23_12 <= vwire_23_12;
		vreg_23_13 <= vwire_23_13;
		vreg_23_14 <= vwire_23_14;
		vreg_23_15 <= vwire_23_15;
		vreg_23_16 <= vwire_23_16;
		vreg_23_17 <= vwire_23_17;
		vreg_23_18 <= vwire_23_18;
		vreg_23_19 <= vwire_23_19;
		vreg_23_20 <= vwire_23_20;
		vreg_23_21 <= vwire_23_21;
		vreg_23_22 <= vwire_23_22;
		vreg_23_23 <= vwire_23_23;
		vreg_23_24 <= vwire_23_24;
		vreg_23_25 <= vwire_23_25;
		vreg_23_26 <= vwire_23_26;
		vreg_23_27 <= vwire_23_27;
		vreg_23_28 <= vwire_23_28;
		vreg_23_29 <= vwire_23_29;
		vreg_23_30 <= vwire_23_30;
		vreg_23_31 <= vwire_23_31;
		vreg_23_32 <= vwire_23_32;
		vreg_23_33 <= vwire_23_33;
		vreg_23_34 <= vwire_23_34;
		vreg_23_35 <= vwire_23_35;
		vreg_23_36 <= vwire_23_36;
		vreg_23_37 <= vwire_23_37;
		vreg_23_38 <= vwire_23_38;
		vreg_23_39 <= vwire_23_39;
		vreg_23_40 <= vwire_23_40;
		vreg_23_41 <= vwire_23_41;
		vreg_23_42 <= vwire_23_42;
		vreg_23_43 <= vwire_23_43;
		vreg_23_44 <= vwire_23_44;
		vreg_23_45 <= vwire_23_45;
		vreg_23_46 <= vwire_23_46;
		vreg_23_47 <= vwire_23_47;
		vreg_23_48 <= vwire_23_48;
		vreg_23_49 <= vwire_23_49;
		vreg_24_0 <= vwire_24_0;
		vreg_24_1 <= vwire_24_1;
		vreg_24_2 <= vwire_24_2;
		vreg_24_3 <= vwire_24_3;
		vreg_24_4 <= vwire_24_4;
		vreg_24_5 <= vwire_24_5;
		vreg_24_6 <= vwire_24_6;
		vreg_24_7 <= vwire_24_7;
		vreg_24_8 <= vwire_24_8;
		vreg_24_9 <= vwire_24_9;
		vreg_24_10 <= vwire_24_10;
		vreg_24_11 <= vwire_24_11;
		vreg_24_12 <= vwire_24_12;
		vreg_24_13 <= vwire_24_13;
		vreg_24_14 <= vwire_24_14;
		vreg_24_15 <= vwire_24_15;
		vreg_24_16 <= vwire_24_16;
		vreg_24_17 <= vwire_24_17;
		vreg_24_18 <= vwire_24_18;
		vreg_24_19 <= vwire_24_19;
		vreg_24_20 <= vwire_24_20;
		vreg_24_21 <= vwire_24_21;
		vreg_24_22 <= vwire_24_22;
		vreg_24_23 <= vwire_24_23;
		vreg_24_24 <= vwire_24_24;
		vreg_24_25 <= vwire_24_25;
		vreg_24_26 <= vwire_24_26;
		vreg_24_27 <= vwire_24_27;
		vreg_24_28 <= vwire_24_28;
		vreg_24_29 <= vwire_24_29;
		vreg_24_30 <= vwire_24_30;
		vreg_24_31 <= vwire_24_31;
		vreg_24_32 <= vwire_24_32;
		vreg_24_33 <= vwire_24_33;
		vreg_24_34 <= vwire_24_34;
		vreg_24_35 <= vwire_24_35;
		vreg_24_36 <= vwire_24_36;
		vreg_24_37 <= vwire_24_37;
		vreg_24_38 <= vwire_24_38;
		vreg_24_39 <= vwire_24_39;
		vreg_24_40 <= vwire_24_40;
		vreg_24_41 <= vwire_24_41;
		vreg_24_42 <= vwire_24_42;
		vreg_24_43 <= vwire_24_43;
		vreg_24_44 <= vwire_24_44;
		vreg_24_45 <= vwire_24_45;
		vreg_24_46 <= vwire_24_46;
		vreg_24_47 <= vwire_24_47;
		vreg_24_48 <= vwire_24_48;
		vreg_24_49 <= vwire_24_49;
		vreg_25_0 <= vwire_25_0;
		vreg_25_1 <= vwire_25_1;
		vreg_25_2 <= vwire_25_2;
		vreg_25_3 <= vwire_25_3;
		vreg_25_4 <= vwire_25_4;
		vreg_25_5 <= vwire_25_5;
		vreg_25_6 <= vwire_25_6;
		vreg_25_7 <= vwire_25_7;
		vreg_25_8 <= vwire_25_8;
		vreg_25_9 <= vwire_25_9;
		vreg_25_10 <= vwire_25_10;
		vreg_25_11 <= vwire_25_11;
		vreg_25_12 <= vwire_25_12;
		vreg_25_13 <= vwire_25_13;
		vreg_25_14 <= vwire_25_14;
		vreg_25_15 <= vwire_25_15;
		vreg_25_16 <= vwire_25_16;
		vreg_25_17 <= vwire_25_17;
		vreg_25_18 <= vwire_25_18;
		vreg_25_19 <= vwire_25_19;
		vreg_25_20 <= vwire_25_20;
		vreg_25_21 <= vwire_25_21;
		vreg_25_22 <= vwire_25_22;
		vreg_25_23 <= vwire_25_23;
		vreg_25_24 <= vwire_25_24;
		vreg_25_25 <= vwire_25_25;
		vreg_25_26 <= vwire_25_26;
		vreg_25_27 <= vwire_25_27;
		vreg_25_28 <= vwire_25_28;
		vreg_25_29 <= vwire_25_29;
		vreg_25_30 <= vwire_25_30;
		vreg_25_31 <= vwire_25_31;
		vreg_25_32 <= vwire_25_32;
		vreg_25_33 <= vwire_25_33;
		vreg_25_34 <= vwire_25_34;
		vreg_25_35 <= vwire_25_35;
		vreg_25_36 <= vwire_25_36;
		vreg_25_37 <= vwire_25_37;
		vreg_25_38 <= vwire_25_38;
		vreg_25_39 <= vwire_25_39;
		vreg_25_40 <= vwire_25_40;
		vreg_25_41 <= vwire_25_41;
		vreg_25_42 <= vwire_25_42;
		vreg_25_43 <= vwire_25_43;
		vreg_25_44 <= vwire_25_44;
		vreg_25_45 <= vwire_25_45;
		vreg_25_46 <= vwire_25_46;
		vreg_25_47 <= vwire_25_47;
		vreg_25_48 <= vwire_25_48;
		vreg_25_49 <= vwire_25_49;
		vreg_26_0 <= vwire_26_0;
		vreg_26_1 <= vwire_26_1;
		vreg_26_2 <= vwire_26_2;
		vreg_26_3 <= vwire_26_3;
		vreg_26_4 <= vwire_26_4;
		vreg_26_5 <= vwire_26_5;
		vreg_26_6 <= vwire_26_6;
		vreg_26_7 <= vwire_26_7;
		vreg_26_8 <= vwire_26_8;
		vreg_26_9 <= vwire_26_9;
		vreg_26_10 <= vwire_26_10;
		vreg_26_11 <= vwire_26_11;
		vreg_26_12 <= vwire_26_12;
		vreg_26_13 <= vwire_26_13;
		vreg_26_14 <= vwire_26_14;
		vreg_26_15 <= vwire_26_15;
		vreg_26_16 <= vwire_26_16;
		vreg_26_17 <= vwire_26_17;
		vreg_26_18 <= vwire_26_18;
		vreg_26_19 <= vwire_26_19;
		vreg_26_20 <= vwire_26_20;
		vreg_26_21 <= vwire_26_21;
		vreg_26_22 <= vwire_26_22;
		vreg_26_23 <= vwire_26_23;
		vreg_26_24 <= vwire_26_24;
		vreg_26_25 <= vwire_26_25;
		vreg_26_26 <= vwire_26_26;
		vreg_26_27 <= vwire_26_27;
		vreg_26_28 <= vwire_26_28;
		vreg_26_29 <= vwire_26_29;
		vreg_26_30 <= vwire_26_30;
		vreg_26_31 <= vwire_26_31;
		vreg_26_32 <= vwire_26_32;
		vreg_26_33 <= vwire_26_33;
		vreg_26_34 <= vwire_26_34;
		vreg_26_35 <= vwire_26_35;
		vreg_26_36 <= vwire_26_36;
		vreg_26_37 <= vwire_26_37;
		vreg_26_38 <= vwire_26_38;
		vreg_26_39 <= vwire_26_39;
		vreg_26_40 <= vwire_26_40;
		vreg_26_41 <= vwire_26_41;
		vreg_26_42 <= vwire_26_42;
		vreg_26_43 <= vwire_26_43;
		vreg_26_44 <= vwire_26_44;
		vreg_26_45 <= vwire_26_45;
		vreg_26_46 <= vwire_26_46;
		vreg_26_47 <= vwire_26_47;
		vreg_26_48 <= vwire_26_48;
		vreg_26_49 <= vwire_26_49;
		vreg_27_0 <= vwire_27_0;
		vreg_27_1 <= vwire_27_1;
		vreg_27_2 <= vwire_27_2;
		vreg_27_3 <= vwire_27_3;
		vreg_27_4 <= vwire_27_4;
		vreg_27_5 <= vwire_27_5;
		vreg_27_6 <= vwire_27_6;
		vreg_27_7 <= vwire_27_7;
		vreg_27_8 <= vwire_27_8;
		vreg_27_9 <= vwire_27_9;
		vreg_27_10 <= vwire_27_10;
		vreg_27_11 <= vwire_27_11;
		vreg_27_12 <= vwire_27_12;
		vreg_27_13 <= vwire_27_13;
		vreg_27_14 <= vwire_27_14;
		vreg_27_15 <= vwire_27_15;
		vreg_27_16 <= vwire_27_16;
		vreg_27_17 <= vwire_27_17;
		vreg_27_18 <= vwire_27_18;
		vreg_27_19 <= vwire_27_19;
		vreg_27_20 <= vwire_27_20;
		vreg_27_21 <= vwire_27_21;
		vreg_27_22 <= vwire_27_22;
		vreg_27_23 <= vwire_27_23;
		vreg_27_24 <= vwire_27_24;
		vreg_27_25 <= vwire_27_25;
		vreg_27_26 <= vwire_27_26;
		vreg_27_27 <= vwire_27_27;
		vreg_27_28 <= vwire_27_28;
		vreg_27_29 <= vwire_27_29;
		vreg_27_30 <= vwire_27_30;
		vreg_27_31 <= vwire_27_31;
		vreg_27_32 <= vwire_27_32;
		vreg_27_33 <= vwire_27_33;
		vreg_27_34 <= vwire_27_34;
		vreg_27_35 <= vwire_27_35;
		vreg_27_36 <= vwire_27_36;
		vreg_27_37 <= vwire_27_37;
		vreg_27_38 <= vwire_27_38;
		vreg_27_39 <= vwire_27_39;
		vreg_27_40 <= vwire_27_40;
		vreg_27_41 <= vwire_27_41;
		vreg_27_42 <= vwire_27_42;
		vreg_27_43 <= vwire_27_43;
		vreg_27_44 <= vwire_27_44;
		vreg_27_45 <= vwire_27_45;
		vreg_27_46 <= vwire_27_46;
		vreg_27_47 <= vwire_27_47;
		vreg_27_48 <= vwire_27_48;
		vreg_27_49 <= vwire_27_49;
		vreg_28_0 <= vwire_28_0;
		vreg_28_1 <= vwire_28_1;
		vreg_28_2 <= vwire_28_2;
		vreg_28_3 <= vwire_28_3;
		vreg_28_4 <= vwire_28_4;
		vreg_28_5 <= vwire_28_5;
		vreg_28_6 <= vwire_28_6;
		vreg_28_7 <= vwire_28_7;
		vreg_28_8 <= vwire_28_8;
		vreg_28_9 <= vwire_28_9;
		vreg_28_10 <= vwire_28_10;
		vreg_28_11 <= vwire_28_11;
		vreg_28_12 <= vwire_28_12;
		vreg_28_13 <= vwire_28_13;
		vreg_28_14 <= vwire_28_14;
		vreg_28_15 <= vwire_28_15;
		vreg_28_16 <= vwire_28_16;
		vreg_28_17 <= vwire_28_17;
		vreg_28_18 <= vwire_28_18;
		vreg_28_19 <= vwire_28_19;
		vreg_28_20 <= vwire_28_20;
		vreg_28_21 <= vwire_28_21;
		vreg_28_22 <= vwire_28_22;
		vreg_28_23 <= vwire_28_23;
		vreg_28_24 <= vwire_28_24;
		vreg_28_25 <= vwire_28_25;
		vreg_28_26 <= vwire_28_26;
		vreg_28_27 <= vwire_28_27;
		vreg_28_28 <= vwire_28_28;
		vreg_28_29 <= vwire_28_29;
		vreg_28_30 <= vwire_28_30;
		vreg_28_31 <= vwire_28_31;
		vreg_28_32 <= vwire_28_32;
		vreg_28_33 <= vwire_28_33;
		vreg_28_34 <= vwire_28_34;
		vreg_28_35 <= vwire_28_35;
		vreg_28_36 <= vwire_28_36;
		vreg_28_37 <= vwire_28_37;
		vreg_28_38 <= vwire_28_38;
		vreg_28_39 <= vwire_28_39;
		vreg_28_40 <= vwire_28_40;
		vreg_28_41 <= vwire_28_41;
		vreg_28_42 <= vwire_28_42;
		vreg_28_43 <= vwire_28_43;
		vreg_28_44 <= vwire_28_44;
		vreg_28_45 <= vwire_28_45;
		vreg_28_46 <= vwire_28_46;
		vreg_28_47 <= vwire_28_47;
		vreg_28_48 <= vwire_28_48;
		vreg_28_49 <= vwire_28_49;
		vreg_29_0 <= vwire_29_0;
		vreg_29_1 <= vwire_29_1;
		vreg_29_2 <= vwire_29_2;
		vreg_29_3 <= vwire_29_3;
		vreg_29_4 <= vwire_29_4;
		vreg_29_5 <= vwire_29_5;
		vreg_29_6 <= vwire_29_6;
		vreg_29_7 <= vwire_29_7;
		vreg_29_8 <= vwire_29_8;
		vreg_29_9 <= vwire_29_9;
		vreg_29_10 <= vwire_29_10;
		vreg_29_11 <= vwire_29_11;
		vreg_29_12 <= vwire_29_12;
		vreg_29_13 <= vwire_29_13;
		vreg_29_14 <= vwire_29_14;
		vreg_29_15 <= vwire_29_15;
		vreg_29_16 <= vwire_29_16;
		vreg_29_17 <= vwire_29_17;
		vreg_29_18 <= vwire_29_18;
		vreg_29_19 <= vwire_29_19;
		vreg_29_20 <= vwire_29_20;
		vreg_29_21 <= vwire_29_21;
		vreg_29_22 <= vwire_29_22;
		vreg_29_23 <= vwire_29_23;
		vreg_29_24 <= vwire_29_24;
		vreg_29_25 <= vwire_29_25;
		vreg_29_26 <= vwire_29_26;
		vreg_29_27 <= vwire_29_27;
		vreg_29_28 <= vwire_29_28;
		vreg_29_29 <= vwire_29_29;
		vreg_29_30 <= vwire_29_30;
		vreg_29_31 <= vwire_29_31;
		vreg_29_32 <= vwire_29_32;
		vreg_29_33 <= vwire_29_33;
		vreg_29_34 <= vwire_29_34;
		vreg_29_35 <= vwire_29_35;
		vreg_29_36 <= vwire_29_36;
		vreg_29_37 <= vwire_29_37;
		vreg_29_38 <= vwire_29_38;
		vreg_29_39 <= vwire_29_39;
		vreg_29_40 <= vwire_29_40;
		vreg_29_41 <= vwire_29_41;
		vreg_29_42 <= vwire_29_42;
		vreg_29_43 <= vwire_29_43;
		vreg_29_44 <= vwire_29_44;
		vreg_29_45 <= vwire_29_45;
		vreg_29_46 <= vwire_29_46;
		vreg_29_47 <= vwire_29_47;
		vreg_29_48 <= vwire_29_48;
		vreg_29_49 <= vwire_29_49;
		vreg_30_0 <= vwire_30_0;
		vreg_30_1 <= vwire_30_1;
		vreg_30_2 <= vwire_30_2;
		vreg_30_3 <= vwire_30_3;
		vreg_30_4 <= vwire_30_4;
		vreg_30_5 <= vwire_30_5;
		vreg_30_6 <= vwire_30_6;
		vreg_30_7 <= vwire_30_7;
		vreg_30_8 <= vwire_30_8;
		vreg_30_9 <= vwire_30_9;
		vreg_30_10 <= vwire_30_10;
		vreg_30_11 <= vwire_30_11;
		vreg_30_12 <= vwire_30_12;
		vreg_30_13 <= vwire_30_13;
		vreg_30_14 <= vwire_30_14;
		vreg_30_15 <= vwire_30_15;
		vreg_30_16 <= vwire_30_16;
		vreg_30_17 <= vwire_30_17;
		vreg_30_18 <= vwire_30_18;
		vreg_30_19 <= vwire_30_19;
		vreg_30_20 <= vwire_30_20;
		vreg_30_21 <= vwire_30_21;
		vreg_30_22 <= vwire_30_22;
		vreg_30_23 <= vwire_30_23;
		vreg_30_24 <= vwire_30_24;
		vreg_30_25 <= vwire_30_25;
		vreg_30_26 <= vwire_30_26;
		vreg_30_27 <= vwire_30_27;
		vreg_30_28 <= vwire_30_28;
		vreg_30_29 <= vwire_30_29;
		vreg_30_30 <= vwire_30_30;
		vreg_30_31 <= vwire_30_31;
		vreg_30_32 <= vwire_30_32;
		vreg_30_33 <= vwire_30_33;
		vreg_30_34 <= vwire_30_34;
		vreg_30_35 <= vwire_30_35;
		vreg_30_36 <= vwire_30_36;
		vreg_30_37 <= vwire_30_37;
		vreg_30_38 <= vwire_30_38;
		vreg_30_39 <= vwire_30_39;
		vreg_30_40 <= vwire_30_40;
		vreg_30_41 <= vwire_30_41;
		vreg_30_42 <= vwire_30_42;
		vreg_30_43 <= vwire_30_43;
		vreg_30_44 <= vwire_30_44;
		vreg_30_45 <= vwire_30_45;
		vreg_30_46 <= vwire_30_46;
		vreg_30_47 <= vwire_30_47;
		vreg_30_48 <= vwire_30_48;
		vreg_30_49 <= vwire_30_49;
		vreg_31_0 <= vwire_31_0;
		vreg_31_1 <= vwire_31_1;
		vreg_31_2 <= vwire_31_2;
		vreg_31_3 <= vwire_31_3;
		vreg_31_4 <= vwire_31_4;
		vreg_31_5 <= vwire_31_5;
		vreg_31_6 <= vwire_31_6;
		vreg_31_7 <= vwire_31_7;
		vreg_31_8 <= vwire_31_8;
		vreg_31_9 <= vwire_31_9;
		vreg_31_10 <= vwire_31_10;
		vreg_31_11 <= vwire_31_11;
		vreg_31_12 <= vwire_31_12;
		vreg_31_13 <= vwire_31_13;
		vreg_31_14 <= vwire_31_14;
		vreg_31_15 <= vwire_31_15;
		vreg_31_16 <= vwire_31_16;
		vreg_31_17 <= vwire_31_17;
		vreg_31_18 <= vwire_31_18;
		vreg_31_19 <= vwire_31_19;
		vreg_31_20 <= vwire_31_20;
		vreg_31_21 <= vwire_31_21;
		vreg_31_22 <= vwire_31_22;
		vreg_31_23 <= vwire_31_23;
		vreg_31_24 <= vwire_31_24;
		vreg_31_25 <= vwire_31_25;
		vreg_31_26 <= vwire_31_26;
		vreg_31_27 <= vwire_31_27;
		vreg_31_28 <= vwire_31_28;
		vreg_31_29 <= vwire_31_29;
		vreg_31_30 <= vwire_31_30;
		vreg_31_31 <= vwire_31_31;
		vreg_31_32 <= vwire_31_32;
		vreg_31_33 <= vwire_31_33;
		vreg_31_34 <= vwire_31_34;
		vreg_31_35 <= vwire_31_35;
		vreg_31_36 <= vwire_31_36;
		vreg_31_37 <= vwire_31_37;
		vreg_31_38 <= vwire_31_38;
		vreg_31_39 <= vwire_31_39;
		vreg_31_40 <= vwire_31_40;
		vreg_31_41 <= vwire_31_41;
		vreg_31_42 <= vwire_31_42;
		vreg_31_43 <= vwire_31_43;
		vreg_31_44 <= vwire_31_44;
		vreg_31_45 <= vwire_31_45;
		vreg_31_46 <= vwire_31_46;
		vreg_31_47 <= vwire_31_47;
		vreg_31_48 <= vwire_31_48;
		vreg_31_49 <= vwire_31_49;
		vreg_32_0 <= vwire_32_0;
		vreg_32_1 <= vwire_32_1;
		vreg_32_2 <= vwire_32_2;
		vreg_32_3 <= vwire_32_3;
		vreg_32_4 <= vwire_32_4;
		vreg_32_5 <= vwire_32_5;
		vreg_32_6 <= vwire_32_6;
		vreg_32_7 <= vwire_32_7;
		vreg_32_8 <= vwire_32_8;
		vreg_32_9 <= vwire_32_9;
		vreg_32_10 <= vwire_32_10;
		vreg_32_11 <= vwire_32_11;
		vreg_32_12 <= vwire_32_12;
		vreg_32_13 <= vwire_32_13;
		vreg_32_14 <= vwire_32_14;
		vreg_32_15 <= vwire_32_15;
		vreg_32_16 <= vwire_32_16;
		vreg_32_17 <= vwire_32_17;
		vreg_32_18 <= vwire_32_18;
		vreg_32_19 <= vwire_32_19;
		vreg_32_20 <= vwire_32_20;
		vreg_32_21 <= vwire_32_21;
		vreg_32_22 <= vwire_32_22;
		vreg_32_23 <= vwire_32_23;
		vreg_32_24 <= vwire_32_24;
		vreg_32_25 <= vwire_32_25;
		vreg_32_26 <= vwire_32_26;
		vreg_32_27 <= vwire_32_27;
		vreg_32_28 <= vwire_32_28;
		vreg_32_29 <= vwire_32_29;
		vreg_32_30 <= vwire_32_30;
		vreg_32_31 <= vwire_32_31;
		vreg_32_32 <= vwire_32_32;
		vreg_32_33 <= vwire_32_33;
		vreg_32_34 <= vwire_32_34;
		vreg_32_35 <= vwire_32_35;
		vreg_32_36 <= vwire_32_36;
		vreg_32_37 <= vwire_32_37;
		vreg_32_38 <= vwire_32_38;
		vreg_32_39 <= vwire_32_39;
		vreg_32_40 <= vwire_32_40;
		vreg_32_41 <= vwire_32_41;
		vreg_32_42 <= vwire_32_42;
		vreg_32_43 <= vwire_32_43;
		vreg_32_44 <= vwire_32_44;
		vreg_32_45 <= vwire_32_45;
		vreg_32_46 <= vwire_32_46;
		vreg_32_47 <= vwire_32_47;
		vreg_32_48 <= vwire_32_48;
		vreg_32_49 <= vwire_32_49;
		vreg_33_0 <= vwire_33_0;
		vreg_33_1 <= vwire_33_1;
		vreg_33_2 <= vwire_33_2;
		vreg_33_3 <= vwire_33_3;
		vreg_33_4 <= vwire_33_4;
		vreg_33_5 <= vwire_33_5;
		vreg_33_6 <= vwire_33_6;
		vreg_33_7 <= vwire_33_7;
		vreg_33_8 <= vwire_33_8;
		vreg_33_9 <= vwire_33_9;
		vreg_33_10 <= vwire_33_10;
		vreg_33_11 <= vwire_33_11;
		vreg_33_12 <= vwire_33_12;
		vreg_33_13 <= vwire_33_13;
		vreg_33_14 <= vwire_33_14;
		vreg_33_15 <= vwire_33_15;
		vreg_33_16 <= vwire_33_16;
		vreg_33_17 <= vwire_33_17;
		vreg_33_18 <= vwire_33_18;
		vreg_33_19 <= vwire_33_19;
		vreg_33_20 <= vwire_33_20;
		vreg_33_21 <= vwire_33_21;
		vreg_33_22 <= vwire_33_22;
		vreg_33_23 <= vwire_33_23;
		vreg_33_24 <= vwire_33_24;
		vreg_33_25 <= vwire_33_25;
		vreg_33_26 <= vwire_33_26;
		vreg_33_27 <= vwire_33_27;
		vreg_33_28 <= vwire_33_28;
		vreg_33_29 <= vwire_33_29;
		vreg_33_30 <= vwire_33_30;
		vreg_33_31 <= vwire_33_31;
		vreg_33_32 <= vwire_33_32;
		vreg_33_33 <= vwire_33_33;
		vreg_33_34 <= vwire_33_34;
		vreg_33_35 <= vwire_33_35;
		vreg_33_36 <= vwire_33_36;
		vreg_33_37 <= vwire_33_37;
		vreg_33_38 <= vwire_33_38;
		vreg_33_39 <= vwire_33_39;
		vreg_33_40 <= vwire_33_40;
		vreg_33_41 <= vwire_33_41;
		vreg_33_42 <= vwire_33_42;
		vreg_33_43 <= vwire_33_43;
		vreg_33_44 <= vwire_33_44;
		vreg_33_45 <= vwire_33_45;
		vreg_33_46 <= vwire_33_46;
		vreg_33_47 <= vwire_33_47;
		vreg_33_48 <= vwire_33_48;
		vreg_33_49 <= vwire_33_49;
		vreg_34_0 <= vwire_34_0;
		vreg_34_1 <= vwire_34_1;
		vreg_34_2 <= vwire_34_2;
		vreg_34_3 <= vwire_34_3;
		vreg_34_4 <= vwire_34_4;
		vreg_34_5 <= vwire_34_5;
		vreg_34_6 <= vwire_34_6;
		vreg_34_7 <= vwire_34_7;
		vreg_34_8 <= vwire_34_8;
		vreg_34_9 <= vwire_34_9;
		vreg_34_10 <= vwire_34_10;
		vreg_34_11 <= vwire_34_11;
		vreg_34_12 <= vwire_34_12;
		vreg_34_13 <= vwire_34_13;
		vreg_34_14 <= vwire_34_14;
		vreg_34_15 <= vwire_34_15;
		vreg_34_16 <= vwire_34_16;
		vreg_34_17 <= vwire_34_17;
		vreg_34_18 <= vwire_34_18;
		vreg_34_19 <= vwire_34_19;
		vreg_34_20 <= vwire_34_20;
		vreg_34_21 <= vwire_34_21;
		vreg_34_22 <= vwire_34_22;
		vreg_34_23 <= vwire_34_23;
		vreg_34_24 <= vwire_34_24;
		vreg_34_25 <= vwire_34_25;
		vreg_34_26 <= vwire_34_26;
		vreg_34_27 <= vwire_34_27;
		vreg_34_28 <= vwire_34_28;
		vreg_34_29 <= vwire_34_29;
		vreg_34_30 <= vwire_34_30;
		vreg_34_31 <= vwire_34_31;
		vreg_34_32 <= vwire_34_32;
		vreg_34_33 <= vwire_34_33;
		vreg_34_34 <= vwire_34_34;
		vreg_34_35 <= vwire_34_35;
		vreg_34_36 <= vwire_34_36;
		vreg_34_37 <= vwire_34_37;
		vreg_34_38 <= vwire_34_38;
		vreg_34_39 <= vwire_34_39;
		vreg_34_40 <= vwire_34_40;
		vreg_34_41 <= vwire_34_41;
		vreg_34_42 <= vwire_34_42;
		vreg_34_43 <= vwire_34_43;
		vreg_34_44 <= vwire_34_44;
		vreg_34_45 <= vwire_34_45;
		vreg_34_46 <= vwire_34_46;
		vreg_34_47 <= vwire_34_47;
		vreg_34_48 <= vwire_34_48;
		vreg_34_49 <= vwire_34_49;
		vreg_35_0 <= vwire_35_0;
		vreg_35_1 <= vwire_35_1;
		vreg_35_2 <= vwire_35_2;
		vreg_35_3 <= vwire_35_3;
		vreg_35_4 <= vwire_35_4;
		vreg_35_5 <= vwire_35_5;
		vreg_35_6 <= vwire_35_6;
		vreg_35_7 <= vwire_35_7;
		vreg_35_8 <= vwire_35_8;
		vreg_35_9 <= vwire_35_9;
		vreg_35_10 <= vwire_35_10;
		vreg_35_11 <= vwire_35_11;
		vreg_35_12 <= vwire_35_12;
		vreg_35_13 <= vwire_35_13;
		vreg_35_14 <= vwire_35_14;
		vreg_35_15 <= vwire_35_15;
		vreg_35_16 <= vwire_35_16;
		vreg_35_17 <= vwire_35_17;
		vreg_35_18 <= vwire_35_18;
		vreg_35_19 <= vwire_35_19;
		vreg_35_20 <= vwire_35_20;
		vreg_35_21 <= vwire_35_21;
		vreg_35_22 <= vwire_35_22;
		vreg_35_23 <= vwire_35_23;
		vreg_35_24 <= vwire_35_24;
		vreg_35_25 <= vwire_35_25;
		vreg_35_26 <= vwire_35_26;
		vreg_35_27 <= vwire_35_27;
		vreg_35_28 <= vwire_35_28;
		vreg_35_29 <= vwire_35_29;
		vreg_35_30 <= vwire_35_30;
		vreg_35_31 <= vwire_35_31;
		vreg_35_32 <= vwire_35_32;
		vreg_35_33 <= vwire_35_33;
		vreg_35_34 <= vwire_35_34;
		vreg_35_35 <= vwire_35_35;
		vreg_35_36 <= vwire_35_36;
		vreg_35_37 <= vwire_35_37;
		vreg_35_38 <= vwire_35_38;
		vreg_35_39 <= vwire_35_39;
		vreg_35_40 <= vwire_35_40;
		vreg_35_41 <= vwire_35_41;
		vreg_35_42 <= vwire_35_42;
		vreg_35_43 <= vwire_35_43;
		vreg_35_44 <= vwire_35_44;
		vreg_35_45 <= vwire_35_45;
		vreg_35_46 <= vwire_35_46;
		vreg_35_47 <= vwire_35_47;
		vreg_35_48 <= vwire_35_48;
		vreg_35_49 <= vwire_35_49;
		vreg_36_0 <= vwire_36_0;
		vreg_36_1 <= vwire_36_1;
		vreg_36_2 <= vwire_36_2;
		vreg_36_3 <= vwire_36_3;
		vreg_36_4 <= vwire_36_4;
		vreg_36_5 <= vwire_36_5;
		vreg_36_6 <= vwire_36_6;
		vreg_36_7 <= vwire_36_7;
		vreg_36_8 <= vwire_36_8;
		vreg_36_9 <= vwire_36_9;
		vreg_36_10 <= vwire_36_10;
		vreg_36_11 <= vwire_36_11;
		vreg_36_12 <= vwire_36_12;
		vreg_36_13 <= vwire_36_13;
		vreg_36_14 <= vwire_36_14;
		vreg_36_15 <= vwire_36_15;
		vreg_36_16 <= vwire_36_16;
		vreg_36_17 <= vwire_36_17;
		vreg_36_18 <= vwire_36_18;
		vreg_36_19 <= vwire_36_19;
		vreg_36_20 <= vwire_36_20;
		vreg_36_21 <= vwire_36_21;
		vreg_36_22 <= vwire_36_22;
		vreg_36_23 <= vwire_36_23;
		vreg_36_24 <= vwire_36_24;
		vreg_36_25 <= vwire_36_25;
		vreg_36_26 <= vwire_36_26;
		vreg_36_27 <= vwire_36_27;
		vreg_36_28 <= vwire_36_28;
		vreg_36_29 <= vwire_36_29;
		vreg_36_30 <= vwire_36_30;
		vreg_36_31 <= vwire_36_31;
		vreg_36_32 <= vwire_36_32;
		vreg_36_33 <= vwire_36_33;
		vreg_36_34 <= vwire_36_34;
		vreg_36_35 <= vwire_36_35;
		vreg_36_36 <= vwire_36_36;
		vreg_36_37 <= vwire_36_37;
		vreg_36_38 <= vwire_36_38;
		vreg_36_39 <= vwire_36_39;
		vreg_36_40 <= vwire_36_40;
		vreg_36_41 <= vwire_36_41;
		vreg_36_42 <= vwire_36_42;
		vreg_36_43 <= vwire_36_43;
		vreg_36_44 <= vwire_36_44;
		vreg_36_45 <= vwire_36_45;
		vreg_36_46 <= vwire_36_46;
		vreg_36_47 <= vwire_36_47;
		vreg_36_48 <= vwire_36_48;
		vreg_36_49 <= vwire_36_49;
		vreg_37_0 <= vwire_37_0;
		vreg_37_1 <= vwire_37_1;
		vreg_37_2 <= vwire_37_2;
		vreg_37_3 <= vwire_37_3;
		vreg_37_4 <= vwire_37_4;
		vreg_37_5 <= vwire_37_5;
		vreg_37_6 <= vwire_37_6;
		vreg_37_7 <= vwire_37_7;
		vreg_37_8 <= vwire_37_8;
		vreg_37_9 <= vwire_37_9;
		vreg_37_10 <= vwire_37_10;
		vreg_37_11 <= vwire_37_11;
		vreg_37_12 <= vwire_37_12;
		vreg_37_13 <= vwire_37_13;
		vreg_37_14 <= vwire_37_14;
		vreg_37_15 <= vwire_37_15;
		vreg_37_16 <= vwire_37_16;
		vreg_37_17 <= vwire_37_17;
		vreg_37_18 <= vwire_37_18;
		vreg_37_19 <= vwire_37_19;
		vreg_37_20 <= vwire_37_20;
		vreg_37_21 <= vwire_37_21;
		vreg_37_22 <= vwire_37_22;
		vreg_37_23 <= vwire_37_23;
		vreg_37_24 <= vwire_37_24;
		vreg_37_25 <= vwire_37_25;
		vreg_37_26 <= vwire_37_26;
		vreg_37_27 <= vwire_37_27;
		vreg_37_28 <= vwire_37_28;
		vreg_37_29 <= vwire_37_29;
		vreg_37_30 <= vwire_37_30;
		vreg_37_31 <= vwire_37_31;
		vreg_37_32 <= vwire_37_32;
		vreg_37_33 <= vwire_37_33;
		vreg_37_34 <= vwire_37_34;
		vreg_37_35 <= vwire_37_35;
		vreg_37_36 <= vwire_37_36;
		vreg_37_37 <= vwire_37_37;
		vreg_37_38 <= vwire_37_38;
		vreg_37_39 <= vwire_37_39;
		vreg_37_40 <= vwire_37_40;
		vreg_37_41 <= vwire_37_41;
		vreg_37_42 <= vwire_37_42;
		vreg_37_43 <= vwire_37_43;
		vreg_37_44 <= vwire_37_44;
		vreg_37_45 <= vwire_37_45;
		vreg_37_46 <= vwire_37_46;
		vreg_37_47 <= vwire_37_47;
		vreg_37_48 <= vwire_37_48;
		vreg_37_49 <= vwire_37_49;
		vreg_38_0 <= vwire_38_0;
		vreg_38_1 <= vwire_38_1;
		vreg_38_2 <= vwire_38_2;
		vreg_38_3 <= vwire_38_3;
		vreg_38_4 <= vwire_38_4;
		vreg_38_5 <= vwire_38_5;
		vreg_38_6 <= vwire_38_6;
		vreg_38_7 <= vwire_38_7;
		vreg_38_8 <= vwire_38_8;
		vreg_38_9 <= vwire_38_9;
		vreg_38_10 <= vwire_38_10;
		vreg_38_11 <= vwire_38_11;
		vreg_38_12 <= vwire_38_12;
		vreg_38_13 <= vwire_38_13;
		vreg_38_14 <= vwire_38_14;
		vreg_38_15 <= vwire_38_15;
		vreg_38_16 <= vwire_38_16;
		vreg_38_17 <= vwire_38_17;
		vreg_38_18 <= vwire_38_18;
		vreg_38_19 <= vwire_38_19;
		vreg_38_20 <= vwire_38_20;
		vreg_38_21 <= vwire_38_21;
		vreg_38_22 <= vwire_38_22;
		vreg_38_23 <= vwire_38_23;
		vreg_38_24 <= vwire_38_24;
		vreg_38_25 <= vwire_38_25;
		vreg_38_26 <= vwire_38_26;
		vreg_38_27 <= vwire_38_27;
		vreg_38_28 <= vwire_38_28;
		vreg_38_29 <= vwire_38_29;
		vreg_38_30 <= vwire_38_30;
		vreg_38_31 <= vwire_38_31;
		vreg_38_32 <= vwire_38_32;
		vreg_38_33 <= vwire_38_33;
		vreg_38_34 <= vwire_38_34;
		vreg_38_35 <= vwire_38_35;
		vreg_38_36 <= vwire_38_36;
		vreg_38_37 <= vwire_38_37;
		vreg_38_38 <= vwire_38_38;
		vreg_38_39 <= vwire_38_39;
		vreg_38_40 <= vwire_38_40;
		vreg_38_41 <= vwire_38_41;
		vreg_38_42 <= vwire_38_42;
		vreg_38_43 <= vwire_38_43;
		vreg_38_44 <= vwire_38_44;
		vreg_38_45 <= vwire_38_45;
		vreg_38_46 <= vwire_38_46;
		vreg_38_47 <= vwire_38_47;
		vreg_38_48 <= vwire_38_48;
		vreg_38_49 <= vwire_38_49;
		vreg_39_0 <= vwire_39_0;
		vreg_39_1 <= vwire_39_1;
		vreg_39_2 <= vwire_39_2;
		vreg_39_3 <= vwire_39_3;
		vreg_39_4 <= vwire_39_4;
		vreg_39_5 <= vwire_39_5;
		vreg_39_6 <= vwire_39_6;
		vreg_39_7 <= vwire_39_7;
		vreg_39_8 <= vwire_39_8;
		vreg_39_9 <= vwire_39_9;
		vreg_39_10 <= vwire_39_10;
		vreg_39_11 <= vwire_39_11;
		vreg_39_12 <= vwire_39_12;
		vreg_39_13 <= vwire_39_13;
		vreg_39_14 <= vwire_39_14;
		vreg_39_15 <= vwire_39_15;
		vreg_39_16 <= vwire_39_16;
		vreg_39_17 <= vwire_39_17;
		vreg_39_18 <= vwire_39_18;
		vreg_39_19 <= vwire_39_19;
		vreg_39_20 <= vwire_39_20;
		vreg_39_21 <= vwire_39_21;
		vreg_39_22 <= vwire_39_22;
		vreg_39_23 <= vwire_39_23;
		vreg_39_24 <= vwire_39_24;
		vreg_39_25 <= vwire_39_25;
		vreg_39_26 <= vwire_39_26;
		vreg_39_27 <= vwire_39_27;
		vreg_39_28 <= vwire_39_28;
		vreg_39_29 <= vwire_39_29;
		vreg_39_30 <= vwire_39_30;
		vreg_39_31 <= vwire_39_31;
		vreg_39_32 <= vwire_39_32;
		vreg_39_33 <= vwire_39_33;
		vreg_39_34 <= vwire_39_34;
		vreg_39_35 <= vwire_39_35;
		vreg_39_36 <= vwire_39_36;
		vreg_39_37 <= vwire_39_37;
		vreg_39_38 <= vwire_39_38;
		vreg_39_39 <= vwire_39_39;
		vreg_39_40 <= vwire_39_40;
		vreg_39_41 <= vwire_39_41;
		vreg_39_42 <= vwire_39_42;
		vreg_39_43 <= vwire_39_43;
		vreg_39_44 <= vwire_39_44;
		vreg_39_45 <= vwire_39_45;
		vreg_39_46 <= vwire_39_46;
		vreg_39_47 <= vwire_39_47;
		vreg_39_48 <= vwire_39_48;
		vreg_39_49 <= vwire_39_49;
		vreg_40_0 <= vwire_40_0;
		vreg_40_1 <= vwire_40_1;
		vreg_40_2 <= vwire_40_2;
		vreg_40_3 <= vwire_40_3;
		vreg_40_4 <= vwire_40_4;
		vreg_40_5 <= vwire_40_5;
		vreg_40_6 <= vwire_40_6;
		vreg_40_7 <= vwire_40_7;
		vreg_40_8 <= vwire_40_8;
		vreg_40_9 <= vwire_40_9;
		vreg_40_10 <= vwire_40_10;
		vreg_40_11 <= vwire_40_11;
		vreg_40_12 <= vwire_40_12;
		vreg_40_13 <= vwire_40_13;
		vreg_40_14 <= vwire_40_14;
		vreg_40_15 <= vwire_40_15;
		vreg_40_16 <= vwire_40_16;
		vreg_40_17 <= vwire_40_17;
		vreg_40_18 <= vwire_40_18;
		vreg_40_19 <= vwire_40_19;
		vreg_40_20 <= vwire_40_20;
		vreg_40_21 <= vwire_40_21;
		vreg_40_22 <= vwire_40_22;
		vreg_40_23 <= vwire_40_23;
		vreg_40_24 <= vwire_40_24;
		vreg_40_25 <= vwire_40_25;
		vreg_40_26 <= vwire_40_26;
		vreg_40_27 <= vwire_40_27;
		vreg_40_28 <= vwire_40_28;
		vreg_40_29 <= vwire_40_29;
		vreg_40_30 <= vwire_40_30;
		vreg_40_31 <= vwire_40_31;
		vreg_40_32 <= vwire_40_32;
		vreg_40_33 <= vwire_40_33;
		vreg_40_34 <= vwire_40_34;
		vreg_40_35 <= vwire_40_35;
		vreg_40_36 <= vwire_40_36;
		vreg_40_37 <= vwire_40_37;
		vreg_40_38 <= vwire_40_38;
		vreg_40_39 <= vwire_40_39;
		vreg_40_40 <= vwire_40_40;
		vreg_40_41 <= vwire_40_41;
		vreg_40_42 <= vwire_40_42;
		vreg_40_43 <= vwire_40_43;
		vreg_40_44 <= vwire_40_44;
		vreg_40_45 <= vwire_40_45;
		vreg_40_46 <= vwire_40_46;
		vreg_40_47 <= vwire_40_47;
		vreg_40_48 <= vwire_40_48;
		vreg_40_49 <= vwire_40_49;
		vreg_41_0 <= vwire_41_0;
		vreg_41_1 <= vwire_41_1;
		vreg_41_2 <= vwire_41_2;
		vreg_41_3 <= vwire_41_3;
		vreg_41_4 <= vwire_41_4;
		vreg_41_5 <= vwire_41_5;
		vreg_41_6 <= vwire_41_6;
		vreg_41_7 <= vwire_41_7;
		vreg_41_8 <= vwire_41_8;
		vreg_41_9 <= vwire_41_9;
		vreg_41_10 <= vwire_41_10;
		vreg_41_11 <= vwire_41_11;
		vreg_41_12 <= vwire_41_12;
		vreg_41_13 <= vwire_41_13;
		vreg_41_14 <= vwire_41_14;
		vreg_41_15 <= vwire_41_15;
		vreg_41_16 <= vwire_41_16;
		vreg_41_17 <= vwire_41_17;
		vreg_41_18 <= vwire_41_18;
		vreg_41_19 <= vwire_41_19;
		vreg_41_20 <= vwire_41_20;
		vreg_41_21 <= vwire_41_21;
		vreg_41_22 <= vwire_41_22;
		vreg_41_23 <= vwire_41_23;
		vreg_41_24 <= vwire_41_24;
		vreg_41_25 <= vwire_41_25;
		vreg_41_26 <= vwire_41_26;
		vreg_41_27 <= vwire_41_27;
		vreg_41_28 <= vwire_41_28;
		vreg_41_29 <= vwire_41_29;
		vreg_41_30 <= vwire_41_30;
		vreg_41_31 <= vwire_41_31;
		vreg_41_32 <= vwire_41_32;
		vreg_41_33 <= vwire_41_33;
		vreg_41_34 <= vwire_41_34;
		vreg_41_35 <= vwire_41_35;
		vreg_41_36 <= vwire_41_36;
		vreg_41_37 <= vwire_41_37;
		vreg_41_38 <= vwire_41_38;
		vreg_41_39 <= vwire_41_39;
		vreg_41_40 <= vwire_41_40;
		vreg_41_41 <= vwire_41_41;
		vreg_41_42 <= vwire_41_42;
		vreg_41_43 <= vwire_41_43;
		vreg_41_44 <= vwire_41_44;
		vreg_41_45 <= vwire_41_45;
		vreg_41_46 <= vwire_41_46;
		vreg_41_47 <= vwire_41_47;
		vreg_41_48 <= vwire_41_48;
		vreg_41_49 <= vwire_41_49;
		vreg_42_0 <= vwire_42_0;
		vreg_42_1 <= vwire_42_1;
		vreg_42_2 <= vwire_42_2;
		vreg_42_3 <= vwire_42_3;
		vreg_42_4 <= vwire_42_4;
		vreg_42_5 <= vwire_42_5;
		vreg_42_6 <= vwire_42_6;
		vreg_42_7 <= vwire_42_7;
		vreg_42_8 <= vwire_42_8;
		vreg_42_9 <= vwire_42_9;
		vreg_42_10 <= vwire_42_10;
		vreg_42_11 <= vwire_42_11;
		vreg_42_12 <= vwire_42_12;
		vreg_42_13 <= vwire_42_13;
		vreg_42_14 <= vwire_42_14;
		vreg_42_15 <= vwire_42_15;
		vreg_42_16 <= vwire_42_16;
		vreg_42_17 <= vwire_42_17;
		vreg_42_18 <= vwire_42_18;
		vreg_42_19 <= vwire_42_19;
		vreg_42_20 <= vwire_42_20;
		vreg_42_21 <= vwire_42_21;
		vreg_42_22 <= vwire_42_22;
		vreg_42_23 <= vwire_42_23;
		vreg_42_24 <= vwire_42_24;
		vreg_42_25 <= vwire_42_25;
		vreg_42_26 <= vwire_42_26;
		vreg_42_27 <= vwire_42_27;
		vreg_42_28 <= vwire_42_28;
		vreg_42_29 <= vwire_42_29;
		vreg_42_30 <= vwire_42_30;
		vreg_42_31 <= vwire_42_31;
		vreg_42_32 <= vwire_42_32;
		vreg_42_33 <= vwire_42_33;
		vreg_42_34 <= vwire_42_34;
		vreg_42_35 <= vwire_42_35;
		vreg_42_36 <= vwire_42_36;
		vreg_42_37 <= vwire_42_37;
		vreg_42_38 <= vwire_42_38;
		vreg_42_39 <= vwire_42_39;
		vreg_42_40 <= vwire_42_40;
		vreg_42_41 <= vwire_42_41;
		vreg_42_42 <= vwire_42_42;
		vreg_42_43 <= vwire_42_43;
		vreg_42_44 <= vwire_42_44;
		vreg_42_45 <= vwire_42_45;
		vreg_42_46 <= vwire_42_46;
		vreg_42_47 <= vwire_42_47;
		vreg_42_48 <= vwire_42_48;
		vreg_42_49 <= vwire_42_49;
		vreg_43_0 <= vwire_43_0;
		vreg_43_1 <= vwire_43_1;
		vreg_43_2 <= vwire_43_2;
		vreg_43_3 <= vwire_43_3;
		vreg_43_4 <= vwire_43_4;
		vreg_43_5 <= vwire_43_5;
		vreg_43_6 <= vwire_43_6;
		vreg_43_7 <= vwire_43_7;
		vreg_43_8 <= vwire_43_8;
		vreg_43_9 <= vwire_43_9;
		vreg_43_10 <= vwire_43_10;
		vreg_43_11 <= vwire_43_11;
		vreg_43_12 <= vwire_43_12;
		vreg_43_13 <= vwire_43_13;
		vreg_43_14 <= vwire_43_14;
		vreg_43_15 <= vwire_43_15;
		vreg_43_16 <= vwire_43_16;
		vreg_43_17 <= vwire_43_17;
		vreg_43_18 <= vwire_43_18;
		vreg_43_19 <= vwire_43_19;
		vreg_43_20 <= vwire_43_20;
		vreg_43_21 <= vwire_43_21;
		vreg_43_22 <= vwire_43_22;
		vreg_43_23 <= vwire_43_23;
		vreg_43_24 <= vwire_43_24;
		vreg_43_25 <= vwire_43_25;
		vreg_43_26 <= vwire_43_26;
		vreg_43_27 <= vwire_43_27;
		vreg_43_28 <= vwire_43_28;
		vreg_43_29 <= vwire_43_29;
		vreg_43_30 <= vwire_43_30;
		vreg_43_31 <= vwire_43_31;
		vreg_43_32 <= vwire_43_32;
		vreg_43_33 <= vwire_43_33;
		vreg_43_34 <= vwire_43_34;
		vreg_43_35 <= vwire_43_35;
		vreg_43_36 <= vwire_43_36;
		vreg_43_37 <= vwire_43_37;
		vreg_43_38 <= vwire_43_38;
		vreg_43_39 <= vwire_43_39;
		vreg_43_40 <= vwire_43_40;
		vreg_43_41 <= vwire_43_41;
		vreg_43_42 <= vwire_43_42;
		vreg_43_43 <= vwire_43_43;
		vreg_43_44 <= vwire_43_44;
		vreg_43_45 <= vwire_43_45;
		vreg_43_46 <= vwire_43_46;
		vreg_43_47 <= vwire_43_47;
		vreg_43_48 <= vwire_43_48;
		vreg_43_49 <= vwire_43_49;
		vreg_44_0 <= vwire_44_0;
		vreg_44_1 <= vwire_44_1;
		vreg_44_2 <= vwire_44_2;
		vreg_44_3 <= vwire_44_3;
		vreg_44_4 <= vwire_44_4;
		vreg_44_5 <= vwire_44_5;
		vreg_44_6 <= vwire_44_6;
		vreg_44_7 <= vwire_44_7;
		vreg_44_8 <= vwire_44_8;
		vreg_44_9 <= vwire_44_9;
		vreg_44_10 <= vwire_44_10;
		vreg_44_11 <= vwire_44_11;
		vreg_44_12 <= vwire_44_12;
		vreg_44_13 <= vwire_44_13;
		vreg_44_14 <= vwire_44_14;
		vreg_44_15 <= vwire_44_15;
		vreg_44_16 <= vwire_44_16;
		vreg_44_17 <= vwire_44_17;
		vreg_44_18 <= vwire_44_18;
		vreg_44_19 <= vwire_44_19;
		vreg_44_20 <= vwire_44_20;
		vreg_44_21 <= vwire_44_21;
		vreg_44_22 <= vwire_44_22;
		vreg_44_23 <= vwire_44_23;
		vreg_44_24 <= vwire_44_24;
		vreg_44_25 <= vwire_44_25;
		vreg_44_26 <= vwire_44_26;
		vreg_44_27 <= vwire_44_27;
		vreg_44_28 <= vwire_44_28;
		vreg_44_29 <= vwire_44_29;
		vreg_44_30 <= vwire_44_30;
		vreg_44_31 <= vwire_44_31;
		vreg_44_32 <= vwire_44_32;
		vreg_44_33 <= vwire_44_33;
		vreg_44_34 <= vwire_44_34;
		vreg_44_35 <= vwire_44_35;
		vreg_44_36 <= vwire_44_36;
		vreg_44_37 <= vwire_44_37;
		vreg_44_38 <= vwire_44_38;
		vreg_44_39 <= vwire_44_39;
		vreg_44_40 <= vwire_44_40;
		vreg_44_41 <= vwire_44_41;
		vreg_44_42 <= vwire_44_42;
		vreg_44_43 <= vwire_44_43;
		vreg_44_44 <= vwire_44_44;
		vreg_44_45 <= vwire_44_45;
		vreg_44_46 <= vwire_44_46;
		vreg_44_47 <= vwire_44_47;
		vreg_44_48 <= vwire_44_48;
		vreg_44_49 <= vwire_44_49;
		vreg_45_0 <= vwire_45_0;
		vreg_45_1 <= vwire_45_1;
		vreg_45_2 <= vwire_45_2;
		vreg_45_3 <= vwire_45_3;
		vreg_45_4 <= vwire_45_4;
		vreg_45_5 <= vwire_45_5;
		vreg_45_6 <= vwire_45_6;
		vreg_45_7 <= vwire_45_7;
		vreg_45_8 <= vwire_45_8;
		vreg_45_9 <= vwire_45_9;
		vreg_45_10 <= vwire_45_10;
		vreg_45_11 <= vwire_45_11;
		vreg_45_12 <= vwire_45_12;
		vreg_45_13 <= vwire_45_13;
		vreg_45_14 <= vwire_45_14;
		vreg_45_15 <= vwire_45_15;
		vreg_45_16 <= vwire_45_16;
		vreg_45_17 <= vwire_45_17;
		vreg_45_18 <= vwire_45_18;
		vreg_45_19 <= vwire_45_19;
		vreg_45_20 <= vwire_45_20;
		vreg_45_21 <= vwire_45_21;
		vreg_45_22 <= vwire_45_22;
		vreg_45_23 <= vwire_45_23;
		vreg_45_24 <= vwire_45_24;
		vreg_45_25 <= vwire_45_25;
		vreg_45_26 <= vwire_45_26;
		vreg_45_27 <= vwire_45_27;
		vreg_45_28 <= vwire_45_28;
		vreg_45_29 <= vwire_45_29;
		vreg_45_30 <= vwire_45_30;
		vreg_45_31 <= vwire_45_31;
		vreg_45_32 <= vwire_45_32;
		vreg_45_33 <= vwire_45_33;
		vreg_45_34 <= vwire_45_34;
		vreg_45_35 <= vwire_45_35;
		vreg_45_36 <= vwire_45_36;
		vreg_45_37 <= vwire_45_37;
		vreg_45_38 <= vwire_45_38;
		vreg_45_39 <= vwire_45_39;
		vreg_45_40 <= vwire_45_40;
		vreg_45_41 <= vwire_45_41;
		vreg_45_42 <= vwire_45_42;
		vreg_45_43 <= vwire_45_43;
		vreg_45_44 <= vwire_45_44;
		vreg_45_45 <= vwire_45_45;
		vreg_45_46 <= vwire_45_46;
		vreg_45_47 <= vwire_45_47;
		vreg_45_48 <= vwire_45_48;
		vreg_45_49 <= vwire_45_49;
		vreg_46_0 <= vwire_46_0;
		vreg_46_1 <= vwire_46_1;
		vreg_46_2 <= vwire_46_2;
		vreg_46_3 <= vwire_46_3;
		vreg_46_4 <= vwire_46_4;
		vreg_46_5 <= vwire_46_5;
		vreg_46_6 <= vwire_46_6;
		vreg_46_7 <= vwire_46_7;
		vreg_46_8 <= vwire_46_8;
		vreg_46_9 <= vwire_46_9;
		vreg_46_10 <= vwire_46_10;
		vreg_46_11 <= vwire_46_11;
		vreg_46_12 <= vwire_46_12;
		vreg_46_13 <= vwire_46_13;
		vreg_46_14 <= vwire_46_14;
		vreg_46_15 <= vwire_46_15;
		vreg_46_16 <= vwire_46_16;
		vreg_46_17 <= vwire_46_17;
		vreg_46_18 <= vwire_46_18;
		vreg_46_19 <= vwire_46_19;
		vreg_46_20 <= vwire_46_20;
		vreg_46_21 <= vwire_46_21;
		vreg_46_22 <= vwire_46_22;
		vreg_46_23 <= vwire_46_23;
		vreg_46_24 <= vwire_46_24;
		vreg_46_25 <= vwire_46_25;
		vreg_46_26 <= vwire_46_26;
		vreg_46_27 <= vwire_46_27;
		vreg_46_28 <= vwire_46_28;
		vreg_46_29 <= vwire_46_29;
		vreg_46_30 <= vwire_46_30;
		vreg_46_31 <= vwire_46_31;
		vreg_46_32 <= vwire_46_32;
		vreg_46_33 <= vwire_46_33;
		vreg_46_34 <= vwire_46_34;
		vreg_46_35 <= vwire_46_35;
		vreg_46_36 <= vwire_46_36;
		vreg_46_37 <= vwire_46_37;
		vreg_46_38 <= vwire_46_38;
		vreg_46_39 <= vwire_46_39;
		vreg_46_40 <= vwire_46_40;
		vreg_46_41 <= vwire_46_41;
		vreg_46_42 <= vwire_46_42;
		vreg_46_43 <= vwire_46_43;
		vreg_46_44 <= vwire_46_44;
		vreg_46_45 <= vwire_46_45;
		vreg_46_46 <= vwire_46_46;
		vreg_46_47 <= vwire_46_47;
		vreg_46_48 <= vwire_46_48;
		vreg_46_49 <= vwire_46_49;
		vreg_47_0 <= vwire_47_0;
		vreg_47_1 <= vwire_47_1;
		vreg_47_2 <= vwire_47_2;
		vreg_47_3 <= vwire_47_3;
		vreg_47_4 <= vwire_47_4;
		vreg_47_5 <= vwire_47_5;
		vreg_47_6 <= vwire_47_6;
		vreg_47_7 <= vwire_47_7;
		vreg_47_8 <= vwire_47_8;
		vreg_47_9 <= vwire_47_9;
		vreg_47_10 <= vwire_47_10;
		vreg_47_11 <= vwire_47_11;
		vreg_47_12 <= vwire_47_12;
		vreg_47_13 <= vwire_47_13;
		vreg_47_14 <= vwire_47_14;
		vreg_47_15 <= vwire_47_15;
		vreg_47_16 <= vwire_47_16;
		vreg_47_17 <= vwire_47_17;
		vreg_47_18 <= vwire_47_18;
		vreg_47_19 <= vwire_47_19;
		vreg_47_20 <= vwire_47_20;
		vreg_47_21 <= vwire_47_21;
		vreg_47_22 <= vwire_47_22;
		vreg_47_23 <= vwire_47_23;
		vreg_47_24 <= vwire_47_24;
		vreg_47_25 <= vwire_47_25;
		vreg_47_26 <= vwire_47_26;
		vreg_47_27 <= vwire_47_27;
		vreg_47_28 <= vwire_47_28;
		vreg_47_29 <= vwire_47_29;
		vreg_47_30 <= vwire_47_30;
		vreg_47_31 <= vwire_47_31;
		vreg_47_32 <= vwire_47_32;
		vreg_47_33 <= vwire_47_33;
		vreg_47_34 <= vwire_47_34;
		vreg_47_35 <= vwire_47_35;
		vreg_47_36 <= vwire_47_36;
		vreg_47_37 <= vwire_47_37;
		vreg_47_38 <= vwire_47_38;
		vreg_47_39 <= vwire_47_39;
		vreg_47_40 <= vwire_47_40;
		vreg_47_41 <= vwire_47_41;
		vreg_47_42 <= vwire_47_42;
		vreg_47_43 <= vwire_47_43;
		vreg_47_44 <= vwire_47_44;
		vreg_47_45 <= vwire_47_45;
		vreg_47_46 <= vwire_47_46;
		vreg_47_47 <= vwire_47_47;
		vreg_47_48 <= vwire_47_48;
		vreg_47_49 <= vwire_47_49;
		vreg_48_0 <= vwire_48_0;
		vreg_48_1 <= vwire_48_1;
		vreg_48_2 <= vwire_48_2;
		vreg_48_3 <= vwire_48_3;
		vreg_48_4 <= vwire_48_4;
		vreg_48_5 <= vwire_48_5;
		vreg_48_6 <= vwire_48_6;
		vreg_48_7 <= vwire_48_7;
		vreg_48_8 <= vwire_48_8;
		vreg_48_9 <= vwire_48_9;
		vreg_48_10 <= vwire_48_10;
		vreg_48_11 <= vwire_48_11;
		vreg_48_12 <= vwire_48_12;
		vreg_48_13 <= vwire_48_13;
		vreg_48_14 <= vwire_48_14;
		vreg_48_15 <= vwire_48_15;
		vreg_48_16 <= vwire_48_16;
		vreg_48_17 <= vwire_48_17;
		vreg_48_18 <= vwire_48_18;
		vreg_48_19 <= vwire_48_19;
		vreg_48_20 <= vwire_48_20;
		vreg_48_21 <= vwire_48_21;
		vreg_48_22 <= vwire_48_22;
		vreg_48_23 <= vwire_48_23;
		vreg_48_24 <= vwire_48_24;
		vreg_48_25 <= vwire_48_25;
		vreg_48_26 <= vwire_48_26;
		vreg_48_27 <= vwire_48_27;
		vreg_48_28 <= vwire_48_28;
		vreg_48_29 <= vwire_48_29;
		vreg_48_30 <= vwire_48_30;
		vreg_48_31 <= vwire_48_31;
		vreg_48_32 <= vwire_48_32;
		vreg_48_33 <= vwire_48_33;
		vreg_48_34 <= vwire_48_34;
		vreg_48_35 <= vwire_48_35;
		vreg_48_36 <= vwire_48_36;
		vreg_48_37 <= vwire_48_37;
		vreg_48_38 <= vwire_48_38;
		vreg_48_39 <= vwire_48_39;
		vreg_48_40 <= vwire_48_40;
		vreg_48_41 <= vwire_48_41;
		vreg_48_42 <= vwire_48_42;
		vreg_48_43 <= vwire_48_43;
		vreg_48_44 <= vwire_48_44;
		vreg_48_45 <= vwire_48_45;
		vreg_48_46 <= vwire_48_46;
		vreg_48_47 <= vwire_48_47;
		vreg_48_48 <= vwire_48_48;
		vreg_48_49 <= vwire_48_49;
		vreg_49_0 <= vwire_49_0;
		vreg_49_1 <= vwire_49_1;
		vreg_49_2 <= vwire_49_2;
		vreg_49_3 <= vwire_49_3;
		vreg_49_4 <= vwire_49_4;
		vreg_49_5 <= vwire_49_5;
		vreg_49_6 <= vwire_49_6;
		vreg_49_7 <= vwire_49_7;
		vreg_49_8 <= vwire_49_8;
		vreg_49_9 <= vwire_49_9;
		vreg_49_10 <= vwire_49_10;
		vreg_49_11 <= vwire_49_11;
		vreg_49_12 <= vwire_49_12;
		vreg_49_13 <= vwire_49_13;
		vreg_49_14 <= vwire_49_14;
		vreg_49_15 <= vwire_49_15;
		vreg_49_16 <= vwire_49_16;
		vreg_49_17 <= vwire_49_17;
		vreg_49_18 <= vwire_49_18;
		vreg_49_19 <= vwire_49_19;
		vreg_49_20 <= vwire_49_20;
		vreg_49_21 <= vwire_49_21;
		vreg_49_22 <= vwire_49_22;
		vreg_49_23 <= vwire_49_23;
		vreg_49_24 <= vwire_49_24;
		vreg_49_25 <= vwire_49_25;
		vreg_49_26 <= vwire_49_26;
		vreg_49_27 <= vwire_49_27;
		vreg_49_28 <= vwire_49_28;
		vreg_49_29 <= vwire_49_29;
		vreg_49_30 <= vwire_49_30;
		vreg_49_31 <= vwire_49_31;
		vreg_49_32 <= vwire_49_32;
		vreg_49_33 <= vwire_49_33;
		vreg_49_34 <= vwire_49_34;
		vreg_49_35 <= vwire_49_35;
		vreg_49_36 <= vwire_49_36;
		vreg_49_37 <= vwire_49_37;
		vreg_49_38 <= vwire_49_38;
		vreg_49_39 <= vwire_49_39;
		vreg_49_40 <= vwire_49_40;
		vreg_49_41 <= vwire_49_41;
		vreg_49_42 <= vwire_49_42;
		vreg_49_43 <= vwire_49_43;
		vreg_49_44 <= vwire_49_44;
		vreg_49_45 <= vwire_49_45;
		vreg_49_46 <= vwire_49_46;
		vreg_49_47 <= vwire_49_47;
		vreg_49_48 <= vwire_49_48;
		vreg_49_49 <= vwire_49_49;
	end

	assign audio_out = vwire_0_0[17:2];
endmodule
