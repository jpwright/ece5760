��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�S����n�Q�<�r0�*[���n��m�"�:���?��Pa��������f�mb�`�T"��f]�����8|m��w</L6��]$�^�$���Bq�7��L/1����hw��S��2�Sm6�h,�a��9�k��ɳ��jz�鸾+��s{��G���aQ7h�w���F<JiU�݁(t��Cw�]x�T�� �0=��VΎS5W��di������sJ�'���^#��i.Ik��(�	����&��׺"�o<)d���*9� �������� 	2�q����=���f���>gmc�ApK�u8�)*e ��<A�$�W�XI���(v螵�wW���j�q�/��`M��1須�ec�T�!�͛� �EA��y���U�d�>�f%���w��Z�	6�-܂ R�����ƽ&Z�t�j���lc��8�/+=���hl��uRe`����f)�q���{�"�����#Y��3?���"%�j��X�������8.l��cTvz��(#�B�(Ƌ"0Q�zb���&�v �t���:$n�մˡ��>&Y{E�>�	=o Y;����45M�+�+`<Eg��o��#�U\�zXS�_�j�0�v��5
�0��	:��i���Zu���*�q?lMa�3u(�{��Z�:��O}�l����g	~����Q��\%�T�Kͩ�j������:��x��5*����t�Q��S���P��0�"��;��Vc(@�*�9�H�ϊ����?��V�%�R���ʺf0Ц�[�|/�5���t!�«�����v���Dm�X�����t GO�^�j%�����쉀>��(�j5��4	k�(\+�0wQ��'�J;c��"���We��ZCK��}HF��s���?��ll�t,j�b�l��/0ܦ��h�g�
<i�ΓpHB1�b��=P�)ܨAop��EO&�~���h7_�м���&�#	��}���]� ~i�{N�O�+{�Kjoj���h2�����Ƈ�uӷ��Rkv��{��8�\J�&�x��@>	�z��Z�E�[�:n���M�٧ ���p���~5D�������֋�=@��� �k��ab���E+�� J1O�wF,=�e�-�P�f��lB��w0�կ���Я�ɕ�=Ք�xg��APtuۭ���Q���p�؍ʂ�.��"�	ihU�y$f}	�\o�NW}������k�,/�(✸�|ʣ�1M�j܀���.[~	S���޿ �z��]����g��x6�TL����<K�;h.D/���8=�1z0ƨ'en�I/4����U����)[d*�`�����DgK� ��D�c%y!���L�v��~�l�w�b�T��6�vu��T�/x=M�k1*6]���8;�$�%����Ko��t�ΒEE��(+�M�h��`&i=R������y�6��v��'s��4:�Cr�$Q�#�x%x��H���������c���D�r����a.��a�7ūF����~�����i�s��h@���Z/&)��̈́	�������O�!+�#��S]m0�֩٘�Z:Ul"�k��6��N!��,=��o�j��!�b"B@H}�x&	����2�B�����A��&�mx�x1����U���"^�&��H�ʔ�<h�BV1�7���&��+ $�s<q�NI��ɇ,�^φ������!'	@Â�%ׄ�M:�!��V����D�"����M���%�ϻ&��3�]B�'[�E  ʃ|�ҋ�a%x1#P�T��]�݅m	Oz[c�����}���2�?���j��`14�0��]ؼ�
������<���%�mឱ�rqP,!��}"��ؾ�Z���+�N/5Ui�8O��;ؕ�v�r-t�h��-�I��@�K�nI�E�TNB�C�dZǕ$ǫ<e�-�h�F5T��3O� paU�j���9�� �V�T����V$�"�z*0������BO ��T �E
��"���!@~�(��@i5����?_+��o�t9�(�=xlx�gX���S� q����]��Gp�A-�4��V}�{���u$����F�J9/��.6�bE��"����u���xڃ�I^�	9�AʾM����V$+�a8�y@|�Tj�����y-���8���e��R�����p�w\U�i�B:k��g�{6r+7��^;�r*��&���/���Q���������V5�f���[K�o��k;��O'9�Υ�ʚ�΅�/��}W��=���oJ���V�sxJ�o��o���<�1�2�yf<�,"�K�(��
�.k�ŐX�N3�
ӓ@�Ww��f���Z�Y������E�*���L2��=�V�|;vYM�8Hv���&ͦ�.y�ͧ*:�l�kj�0���a����
G���@��
l�
�+�'�����|�H��2w��I��kT���R/(�Z�p{��ak
.��]�}�ϔ�f���H:���=/
�b~2��'RY+	*.� k�]��%�yw�8i�3]�Y��$h�rF��Ћ���~�j��P�:]f���@iSӣ����\��t�|��EN��XH�$tC�� ٢������Y|pb�9ho�f7����Ǎ�k�c���(��nP��CbC�ߦ��BQxEKɉ�q�v,\>���'��7f?�ODŵ�;�D���w9^��5�1�������[�w� ��ߪ�MH�x;?f��Lh�������؛���Sa�7�gY/����pS��ߔ��)(3W�]��Y�ε��c�����/t�� x/�6��tE���7ׄ�zW7P��tԻ*< ���33��G/%��Co�*;�oMN���������{�̊��- G�@J8�i��@��}W;��K@��[�c^_��h�|�"M���>{�Hp��P0#+�fm�⵱�i�c�8>�ހ�A�<��0�͆���IW����2Ő���~4��W�0�k�$5-�񻧥��b#�-Z�+��40tT+����Z\��8��u����{#�m%�@���h|�"s%����h�C���+A�i��Vp��<6��a�:�M�t�.��C`f!�8_\��3j�ŧ�x��/�T�^Z�n�$9��_3X�D����z^C��2�a�=���V>�f|��z�+ ���AYg�cp�eD�o�����M���T�d���d���o
7�cu�p���A@�A�'�b@xgơ0����Ut#�9�¢ޡt�P^��i]~���F��`P�g��%��Զ�a�S���)}]�d6| ����e )����t�fq�.��!��Mq߈1�M�$���)�y��vb�,� \�0�N�~C�EE"�v7��!���bj��y�l��T�%?j�~z�y�O8����-z�*��rn�@gmf������\�p�r�4*��61>G�u���z���cyh��sxpGC5&`e���T�U�9��H��.��c�,����~"Guk,d��.�N��ab0<|���U1�9�^�պ�ZZc�Q�Ie ��t��Z� W+�G<I�]�0�zAvv:Đ�3��z�~~<�-�C�;�uc�F���C<�qAv^����Si�tU�!�C=�Vj��@�CX���y&��;��fd�fG�Ġ�AU��ٻ���k���+u�	*K���o1K.��n�Z�,�@���#A� ú��Ԍ�8�u��oʂ��w�f�� �u@����B�hG�؆�S�*Y���m�}�2��_�aJI����Ƹ��!� �bqc!',�D�C컌W��$2W��8"1h�%��'WX��SU�,� /g�z�?*k0R�uJ����x�E07J6�b�A�?�(�Tx�Խ��cVA�)�\���rP�;���3�s���Y��f��p��� kW��\��]��/B�:��~�W�J1�m���
�a����4K��Mp�Si�iP���B�c���{.��Gם�{��tgg��.lLP?#<PL͎�mqc(9�0�n�ߧ�x��gZ.T%��P��{�La���vx�a,cK��f�ou(x���ASZ��8�R^���W1�\�=��_�����ߓ��'�3�ڎY�ٝa��Ι̻3=	�ˠN�cI��?#�&�P�nh������(	�����V1]� �/Y�@�A鹈P4��81϶�0a��(I� ]��t�C2�YL%�Kr��m�Uiǹ�� �M���Nl��`׊:I�_ϡ}���r�"��<�ñ$i^y���G]��Ï�	��	Q�UA	n���l�4}6���t��g%:�<>l_���a-�N� P'�q�6LU��%�]��>�x)�"�M�Q��X4��ӵ-�����lȽ��'������n�]xU]m�L���B��R�^�Ձ��7/��I�\����6*�$�#�$�׉��$�/�M��+-*y8���TU���9j\W��2p@j��#�膔�Od�|��a�!����	Vu]dĳ���YWpc0`;�领12��d޾CF_�X�_¦�x�`�5�{��(�d�ˏ�,f�WK�S�ցFW[ɐ�{�Ӯ�6�KɅR]��;��U��Qm}�U����l�n)-R6i�r@6x��j*�?+�y`���Z>�N�~�����bF�\�p�!an栠yǌ8�-�� ,�+�Ϯ��^ �3QkLi�u��f��`lp��]8Z*j��:�=9�����.$�R��J���rc���h��A���?}x�#Y�����vw��tq����[hl	̙d��;s���,[g֗�`S|&�}�H!�J7�d��]7#�o�V�g|q�Ғ,qk��On�6[�6Sk��m{�DQ�
�և�K{'���})ᰃj2LY�MlAH׏e��J��C	^��0`Ч����HW6��G��"HC[�������*�EgEͰ���<<0邺��F'w�s(��`t0Fצs�'<��t�K�bT���	2#|���I./�q�E���oZm#��j���\�����	=2�F�u�̙ʸSXlu[d m�{S��:�٪�c{܋���RW�^�:��3���X04_
�J�B��89o�l�>������h���{�ս�U��aҋ=,��i���Iyp)5�
v-�{�⥐s�ɳm4��9e�+�4r�R?��$K�k{)�[&���e��|�ɰ�jHw�Q����� Ĭ&�+މIc�$"��$<��C��ejċ�.4�_Ѹܼ{���\�<R[#n��ikV�|])���H���W8���+_LH�7�|0�Y�aT�24�A2^�l����>���c'Q�wS(�K�	����CD�pGV�H/�EH��Ne�n�ȵm���@�K��G��)�h�o�B�X��m�Ƽ�n���y�~M1�����j��e8��b�^�l��7N���{�8��3�2ߗ'���;�檬@���Vp&.��&��L�K��P�Q͸�/����F�r�7ns�L���Tŉ�r��6�[�]sҝm`������� �|�f�s͟�C�(��-bÔ~�4>�SN;�p�͡�X������G��X)�vP ?R?�c�Џ��AIy��q�>�س�/��YB��j��(�+h�N�������}��^ `�ykO������lJ�򟰘 ��r@�o+Ti����76a�Hݺ"!�����xM=�Xة���@Ш�����I���l.G_�ug�ֱ�	p����E���Gn����rj�_l��)yo>$8�W��XY^���'����/�of�5�bo�<c�H�RV�z��=�v�1#l�>���^�W�8�"�"ȶ_T�	!�<���N'�~y� �Z��6;�u�p�}�,8�V�Cᙒ�^oh�9��E3�юS��2?�R��|���*�c�܍G�]�u�$��Cq?b�-��@UYo����ؕ�<����'���}��`h`�ҽ���k�E&a��+�e$:��Ϫ���������;k�[��Ŝ�"��Ui3��梪���h����kH&�����i�!t6T���
�y^a����<�az��=�t�##@'s�1�o /�^ȣ���5��Q�Ibg��[�Ǡ��g�b��������A/���ZۗG���"K��������myJ������=s������v<s��OV���u�ϻ�^��yB<�1���9�~F��N";��=F�ߛ�v��J���ϡ�R��;�hTMk��� �oNg����S�r/PD��Ɣ��uF�Ju���:���+[�s�6��6���/��^���\S�-�+�+B+Y��Ր���B�S��W�n��FK]��1�a���]�Ld"V�z�l�l����t�������4fDQp������Գ�|sQuc�K\F�yk����<d4�=�>�"�S�����ʓ�0�+w�$���ɮ���A�8�A!mR��]����IC���أ�� �cl�;(�!N�t �4��h=
���a�p�Gu&(>��ʲ�4�2ڏ QF>��{D��1�q	b�n�w���5P	'>�j�����-ޣJ�v�a)l2w@�y�T8NN_s��_,b9�NH�ۚUr2v����^4�n��%Ur��-�#eJO4rS�,3�Ebk�r:���� `Ò���g�	N#<BgT�t �! �n!YX*�<�fI�TT��WK4���N�)L��ؼ$H�y��ǣ@�&��)��>���<��sW���AШ�#ARX�% �yi�ݐ�st.��%ߕ5|�B��u��6-a�#��ss0\\^J��6��aq�L�Tڰ�m�i�E�f�uxi��K���>Ɗ��:��g'��F��,� n���K�2f��r8��S;�=͇����뀇�6��~ ��$70|�K�� |�t|�S�DӍ��T��_u�]��)>ql~ ���˴�ltY#/x�=���s�1��ޞޙ6D8�u-=�(���:|Y��k=�"��t�逻>Ͻ�h7��`'h
���֔j�<2m��h �YߛRp+t��@>({�8V����iFz9�!R�Q �R��6�bȼ_����&��'֊?��nY4��@U�����?�����o�2��8�U���j������+�a��>�RF`�I,�7�5Qۣ�{wR�#}��yu��@��B�u��+Y�?���XI)���֒>��Ѥ��YZR}��1�%�0�TR�@oz����H�U����Gb��2�܄�xX��g�����C�^_��?]C�N1B0k�6AT_���d�O��D�V��D~M�޷�)���@��J�7J�&k���UI_!�g��)��o�������ǜ��B2y�ӧ
K�P�&���8�G���O���-2����w��0d���^�4�?(������̡"b����t��T<P%�ċ&b>�M����c�s��(�8J��.5�EH�a��~g�]'F(���T� $ӳ(ˠ@CW���}[�GӢ��]�CN���EG))���>���q����PB8� 8�� �:$	�S)S�,aE%��,�`�F!>m4�YŖY��O��CMk���7��Ʋ�H��
`+H���>� �x��љV�:��Q�!����� PC^R��s3,����9p�9���n>�#e�0"�&}@�7t㢡���*�`k,O���z�y�z�C�,#���eNTD����:���f�9�K��>��e����Ke��㩢�V��_�l�J��l=6�0����i�ZT62^
�;�f�tÂ$��1�[�g)��jn�FM��W�/D�I7��Ҭ="qW%Ehl��z�U_�Im��8�[y4H�������`�H!(���<)��Z�*A���H�[RV�ʞ+���d(�n��������'�v��?j$b�Gτz.�50 ���.�%f۽,B6�N4���7��E��}ݤ��T�)�]�>g��k�R	�oT���
�j�ԃ5U?���u�Tv�;���j�"&n�\Cx���u��@���U؉_�ґ0�l�]����搄�s#:L��ne��qi��\�]��b���5�����O��G�Q��I���o��}y�MH�&8VYB�K�^pw	�X���,�����$K܈j�(�hȨK��d^�S���N�j�~�.H��X�ڞ������3�i:���a~ ���/���6�6�^s�J!j�����-ƅ�a��׷���D��O�z���9�������{�7�(՚��i+�Aw�J�
u�E@B򯥅tӏc�����kN�xaiEGZ�q~�q����V�Q,ƙ��9��{�0��\�/���E���r 
�3G�lC2��ZcЛ��ϊD�X��1k#���@	Uo�e4��%te,X^�t}��w���b��g�?e�KϬk�V�RwC�{��-2����+-7��B���{<���(3��%�4S5�!54)�^M�.���M\ڃ�d�a?���)JK��z��='�th.O7���G���Ϫ2%���j��P�n�<
��7�V���G���N˃{j�2�O�F�b`(�u����L��w�����e�g���jp\v(�Q��	1P�����{ƪj�	tQA�xw���f��[a���2$����vrӌ2���c0ZM�K�zE�@��������6������1�x���}���>���G`P�	�n)�*�nn��K�[z�к�𰇷@�g5�����7��h��,;[s.�A1��	.�D�]��2��W�c���u��dj�LE@�^������?`-«ݨqdғN��Ț�&�٤By�<�GM�ǫXx�8��� �N3b�7�G�ɜO��o����KHrd��|,ZXEƹ��FoK׎���=r�+�M]�n��u^���5j*zh��`�^6���y�9��ccDS���T��k�Ŵ�.���Ps�G[,���ȓ9��J�~Σ�A��Ԛ�c@6[��ƹ�H	��4h#3�jK(�4p]�	���)�R��C�gZ4�d.�3�Y��aߊ6���?��IB��q��j�3`�"&�/j7P��9�=�@a���	0�ІK�+J+�@����L��a���ʦyJ m�-��#"��vi;�Fz�I���}�*k\_i���g2xg���2�b���B:y#��1q^a$��ؚ�
�7])�.��1!�J���6l�_Z[����+��������b��IKҔ�8��*��L�;dDva~ڸ|N[�{iV�F]�}'G"��ײ��N	�%�,g�I�;`�aC��O2�$�9�%:� �M�4��nWPB_��7�)����&������R6����E�𲿇X�>�w���v.�F��PSN�tAyKU�s5�=coyOr�g� ��5Z"����5�C�����OR�`��5p���f@z�������bh�\��C��%�ܢ�8���!��S���ł�z���U#���\ ①���^v�s�@���	�������FV0�O�
��5�h}>A��;I��������xG��`�V������-q��x"�G?��mE�7���ԁ_8�-F�$���V5�E��g��vUefǒ�+���[���ٛ�$�_�[�%��`�p3���t���׸����ml����eo=���2�\�k
��BLj������U9�]\;2w�����T�f�2���1�~�tn�V.~M,�4c�w���d1
����x�TO O�q��>4.�ϳ��������8J��h���M1c�SA�o��dO:�inh�w�P]KX��L����I­�Qj�&��]}�m�{�|��Ս ^��m�V�|��3����@�Qr�р:��n�)��۾��>����]�/Ǆ�F��ξϻ8<<B��>'���dx�����Z9�Fa��1�{TQ�}�F�#_�m�e9����~�����$��q--��O5��z��E�n��*�ŕn)��I�2ߐ�yJ���Kz��RBbu�o#_��YTE	Q&� W��.�乑��s�"??�G.�9K82K�����!	B�%�
����Ss��xY<Yn;�$������{ggJ+����+X %N�z�i����C�+����^+�I���sW$`�1�>~9,|�j�)��?Fq>ō-�@�%�^�Y����0�L��N�T�YN������!��)SFVM���P"�|w]�)��r�=δ�pBCҸ�N��Ä��@6w�\�1�b&��i��8b,e��
1�z�$�Ʊ�V��^y*���-^qWީ��T~Og4�?Y���lo춤���af���T�ٙnC�r�o�P��7ź�������t��k�
RQ����	�6���rȝ��$=kF�R�����l��T7I�c���i�������0�B��p���T�Oՠ���8>}���1R�j<1�J�e+U��;wv�T�5��&"�jI��W�|�{�#X��H]���=z�I�D�\ ��YY���KV�T��'�*�����@�d曞����+ݧY �d|���#w/�v��-z�1��L���,��U�Eg� ,���:���Ѷ�`9\�����N9G����yZQ*W��G���5�i����_D&�Z4]���T��Ѳ��j��LD��lz�u�e���vD�h:� Л����k��V����Pu�d����QL�8c�4O�?A� b������Yw�:�]i�}S�}*�=���M�p[������q��}rp�QBC]�� 1x��A4�bA`���"g�a��M�{2ez�K-)m_�=O��S�Y��������aH��,�:?f�C�'+ϧ�Zf�#���G/�qōx{?�<���@����:�ê(V��I���ҫ|�<�Y��%:bj�_s8D�iZ�
n�|"��o.+�P$2��4QfH�0�El���Ĳ���v
���i;�m}k��1�Sl��E��q��S-�G"���y=`���4��D\�����E���l���Uv��x�q'*��{ˀ�����*��m�i)�A!�	"��5�g����h�FV�9�}4�LX·l� ��o���'Gl3�S'ȓ�����p\�E�0���od��/�Vh��L��"�)��XM��5�U�Z�`WWˀ&��J��D�gh�W2d�q��}�����f 9��W�R���i�(�Ĺ������*.�x�&y�"���W]��ǙD:O&	��K�u�;�(3_� �T'b5��#�M��lߢ�)j��Y��a-a%��T���)]�eĔ0�h.I?�
�R�*��۔5Y{.�$q�-�T}��ȅ4��&�V�1��O�,$�t��b0�u�U�X��d�@�B�&� Q�oq��@ȸ����5� >�w�Ɣp���PF)��,��m_�r^2���N`�+����,"��h��a��ǰ�	��α-�#���s%���r��u�^��y�Zֆ��
���z�x�)��Z�����C��&�)?��"��&&��iZ�b�	|����3���p�����B��{��+�����VC�R��"�/����5���a�
jE���c�W��т,5�����VVa�#6H���L��G\����/�
WY�h���#��:�+�R��0V��1�},��۳#�� CL
��ڤX� P9na���bb�]׺s
x�;� жcݳ�S��N�k;��;K�R�읗�"�x�˙�zδ��ۊCRc�|�=��C9���U�<^U.����	�>����k皇lwy����6���Wbi����,�K1�gy;'��J�T���I��)U�q%7� g����;O�kQ_�-�@�V���.�������}���`v����"4��^�3{�������I �A�wݓ!w�w�V/������+K��#�@����e�f�d
�8��A7�Y@ܖ��k���u���&7��\3��g�m7*�r��[�EJh9F�����xS�Q\��~}��puFY�Yk'�J1i>�� '�5N�� ���v4��[�W�y��Ϥ{ȉ<Sx_�>�����}%�G�i�V�jڱ���+�N�y��G9�E�\:�Q<��߳�\S�7�E�ub��-�`����V�a�v�{��Km�]������0U9����$�!}�Z�����X+��h�n�>�A�O�[� ��<��U���\�`��j�)��{�Al,M�E�`��Q2��c�� �b~\�5*�'���o�c�J)��k��Hꊬ�bHo���,�p��G/���=��np���{���,ՖZ�AU6۹���/�5�����,2��I)�
���|_���1�&�� �#�ᦝ�Q�2�l�
��JhOr{�����U⓴����#Lmp�:��mbO��:	����@B��¿�X':��oz�j�{7iF�Ni�uЦP�%�vzi�I�_f]a���֨�tN��7b	����/Bװ~A�'�J��	���JUG "��X5���bopI>RҸ=�^S�D�F��{��}##ŃB���/hm/����PȕOe�aw Q�к�:��5%ZO�H): F̍o+&Is� ���i	�I���ni'�$o^Xz���}���3���U+@n��G>��=�XvVC��jg�]��sC��L�r>bF�V��NT�<����&�SE�k���C�z ��_���̢s���}�X�ʎ��94���^L{����6�Cʛ��^»`�,4eh?B(���i:�G�-]�-�$ȍ�5C�Jf�Pń��j3�w߭1^0
��ǅ�GR�lV�Rռ5=k� ��Ϭ��Pw�$�h��&'A�VY6�c�� �E��o��4#�||4����n�����U[F<�{��XA4�W�1��mURX��c�r�������fHuz��=���C��a�'Oߠ��\n�.��6���?B��͇I�)�o�F��a���@R���v6��x�y8��,�#���W`�&ǈ���7��)v궨��&>�<�����A>f�{�X^Ԉ'Ԯ>w��aE3���s0�ӎ���'f�B&W���hm~Q�S����'�s��5`{B�:�rLӥ����A��%d���kl��(&^�W8��	�R����'\��)M��|�j�T���r!D�oy�=y�2�Ow�n�l�T�u%9λ[d$��z�p��U�4y[�Uk��]�$U�hœ(�"]#HU��q�����ʓ �	��)1��oF�;,�ŕ|{T����G�P� ]�=05s�2�j.����o��J�=��U51�!�T�:*|�
���^�vҚRB��� �0 p�ks0}L�ֲ].��1X�����)nV�em��G�T�9u,b�u��SH>������,j	Ƥd�;r��r0B0	�A��RB�����gt������;�W��̓]G��<��H�d�VW�;u��ޏU@")�O����E=����v0�^SL7��ͯ'��ԅ��H?z ��R�N��G_]'��)��"�)C�,��=>��$�D%�D�RX��Fӝ������G��wf�,�fW�-�������������t�Ǜ?�ݐ'�ȣ�<Wi�B%3���7�k�Ɓ�Ļ��w����m�ɭ[���������)��r��p����g ���z�T2�u1-����f6��Z�$��_~�Jd�%��՞S��)�a����?&S3����A������'h��(=�щ���S���В8s����D}\ge�NpA���/0ӝغ_���L=��l�-ԕ�l6��G1���2}j'��8��rEy�σ�Qa��{�@Guba��o���E��y�d���E��lw(i�u(����A.�:�A:%�⒔�usq(`t�\'���=Lg3.9s�zN��g�f�.#��3~�)�X�'NE+��ׂ/��X��Q��}PP��?2"��.]��A�M<{'�U�&'1�Ѧ�}�/Un�W�����������C�3�M+:C�xJ�nz��
9����������L��qf�7�K�&,����^�q�9غ�`�q��B��r�܆��ʢm�9_�p)�h�^���
,Ue�6��T�%�9������O���6�)���}�j�@E�F�ҟ��E���`����.�g��R�I�V�sQ&�Ч��G��â1�8�$;m�4�7L��pP]���cP[|w`ꋨ5C5��no���$SMtR�-W��v��x~qWݞ{�,?&uʑ,W(k
P��A��uv��a��)4�HpsmK��6�W���b�������
�����~��%J�/��g2�)6��V¦a�:7jǁ�����j�j����KB�o��3��3�*,�W^~�z7��u����/V��}� ����Z�S]aڥ[������{D�ѓ�*����%�����x�ƭ��rs񻎳��Y�j(�$E��qp
հ��r�
�K*=�؁M���Ct�`x6n����~�����i�+�����o�K��(-j0������Uo�v/�=5��j!��۳M���T8�>�W�
��:­v�9g��{gv�@P�{�A�Κ#x� +�<�ڳp��Յ���o�{����E�.���s��m��MPdTU�gLF1h��b.5a�Y�]����0)`�vհ��A�X7)bű���*1"���z�%QIh��cR;F��N�W��1�М$���JZM:�1_N�J�6���R��*�D�%�`LX�.��yސ������s:�u
�5����VCg8 �g�)���hգ�T%Ʌ��m��jm���e��Ztb6G4����a� R��Y=4���Y*��H� ٭�eSS��M��]C���5,K�7���uh	/J<����}��
M ��F�~�?k�1�QTLY�+��3�]����8�1
E���Aj���:��(�t�*�o���R�����z�#>a�̿e1ߞ�����lu���b�P���9�:�w�)W:�ZВ"Yoi����N@J�s�g�N�;�W	|������{�"Qf�G��_�>��Ra�Fʚ���T�a��(C�;�]�cM�����T��|]Rn�3�x�h�vx\� �d�E���[o}���O�[�S�k���fg�/o�q:�<�9��&�VT�]^17��B�	�Q e����uŁ���бv/\ �i�X!�i�LUI����w"�7�trOZ��d�S�K��i�P��Ef=@�`f�I�P��d���f,&]5���>��~ƞt�3o0��DꐌT(�>4E�t��d���+�j�Յt��-{ /[ �uG�{GI��V�`�����T&!185%5~����۴C������y$���x�z�vӳߐ���Z���n� V���fD=�o���d޵�_	�gm�,i��	).қ�# MI����Ʋ4��a�����,� ~Xj��|ƕ�"fC�g4��`F�M�^���L>�j�y�!t�l�;�W�_:�x�&��J:(ᕚ�vE����þ�d��z��ժ>C��ɵ�~���7-��X�Cs�Y���������k���Y­I���ȀA���2�4��8�Q���xF�%<�O<��l��ߘҞ~�1�a��j��� �b�=����UbC�K�A@~��o�]D;�x��re���t�Jэ7��zA[q���1P)AZ�
����Q�;����Lb˄"I�"��f��q!��x�}�6epl�2��'�٥�Į���>(����=�~�h��
Ad���@R����,��Ok�����.�of�c�Ì7�z뤬�P+z��ew���`�-�x��h��85tMA��[�F�K%O��dI[�7�.�h�	��2�hD­����}�οB��Jߩi��(
H��/KS����-���AM�@;�^�EE�r����aR�J	^N��Ƃ��@"t�*+�y;�B�0��d�)�c%��X)��_�}������B�&�,���xߓ2���Ɲ���������i@E���VX��.YX���'�WF�������c1L���$f�h��$�}[�(����BS�ٽ!u�R/�ﯦ��,�G�cb�2ƛ<w5Co��R�q)_�Đ�CK4�P\Y��&L���kt)S�YB�x��Q��+�Y]�E����]�Zr��@�����a%���@�]L|9�pGMbƒ����<0��=fz��1�s���s��)|Xe�9LW�y�L�] >�Fy%�l����w|]��P�����~&� K������0�z�&f�Lׯ���q�����/�e���ɷ�m��H���-./k|"�^*���M���?:&�� �T���;M$Z��r�?G�>��ѳ%98���`Z�Fd��z�8����p��+D�7;<�9(����:D��8.29��6��9o����>;uJ+�{�Nṗ��%2m�sW�z4�&��_��b�z}6xlo����G A:M�������/d	��m��D�z7�3��Φǻ��/��$8�wTY�b
!�5g�P�����*F��՝�~�����ڠ4詐�y1K��܆��NB��6Ͽ��L����Ha���F�2��nSѰr��� AU��#s��čc�9b�ee-��0��x�Sku����0���ӄ���C��+a�qK�'�CgA�ީ`����?���I����E�~�Q�Fto�r}�ѲR0H��c���vf��S�	�������uu%H�5�rz�.�7e�����3;�>|�F�V{�mC�ϓn��@q��8-*K��J������b����R�����o��PXWӶ�D���KFu�s���"�{f�m�Q��@� �#�v3��P�.�����?�E5��z�Y��@��K�E�"�|�%=C#I��e�3���<�x�䕴�
;��ْG�E�s:߹�� E������^=��H�f�Y��k�L%�(^�SP�)p:��l	� �����W
�B^MKצ�6�Q�U��Jq�+/#���d�m�������όa�5-��3�L�W���D�i	�hB�k�K�G�K)E<a�e�1�Wwg߱ޒ}v@H.6��˷O��(���ȷfs��	��9�K�ԯ���]�f�YEE}"������j���Bw��Ɵ�������l�_%!4�@�
Di�U�	��r�t���\%y9*2����`���T��u����GHZ������,��¨ �9�D�|f�ԛ�S��̙Zku#����8�|��UP�r���YS�vxb@��-�%l���e��|l%�i��Q����/
�qu����]�r���[�U�4J�pK�����"<{Z���F-L�)�΢Au`-\�)�Q���Ұ�KŊ��� c�������Yɍ�t�L4���R̅�cDCAS��x�kJԙ�₩6�n;�=���^8�cJ���;�_jbl4p�j|SY�IG4��̓�4Tf&Ι&PB���֠v&������jV,�$����K�����(Z4�L9��J�F���4C������g92I�5ß��%M�<��a�[�	�5�5_�2��+.��0�bN��gL+�%��$�2Z*��|��C}ȂӪP>g����;p�k����%���6��D��K)V����wz%�K�Aq�;r�Ȼ�����!���Tr�J� 3�kv@e�V6��%����� ���~Z����jh3ZW�|O�"� 1(��Y�Ksߺ��}�� a(��2���u&Mjg
[�g�-k1��1����R}{=��Fho�]J�&>UY�os����UJ�6�S�� х��'�a&{�G���80eʷ�/1U�S��65h�M~7gUVɥ�݌R¶ޔd�x�9n��������^眯�6"��xrە��R{y|.�ׇR�y5�����?��#�6����Q��F�c��Q����*�[0���z�c�V
"*�,l����y�q��\� ��1�Ve�>�]	`)m'wN��1�m�ޥ�w[�P��x�qYzz1�z� ��/�V��~�ZqKB��P80 ��O��!�ҵ�s唃K��1����G��S`8lD�`\P���`����U�I���$��lP����Z����X�6��8�ޠZ��֟yV��'����s�X��.5#\���NϩMM/�=BK�G0ᖉ��t������nd��\>#w{��*�#)x�� c���ʖ����8�Z[�u��AQa������ִ�)�#b�$ �1{b�bC#F>�ޜ�@1��D�^K�ѷk[�F�/���zÌ�@��,>�/+t��dB{��E������O��yP�� ����q���<Y�"����(&���}M��z��i7��o@o�f����9�|��&�E��<TP�0�o�=�2����:�TW���~���OP�h0���o?r�nx>����[��:����*݁�!bC��;��>�Y�"�6�ot���ॲH�D�N���P�y\��Gw�g�A���0�	˰�3�d<{�zU|�\�$�,��r1�}v�������ܳ߿%~�jG��MFf��U��]��E��Q� /C��\���5�+��n/���&M;l׳u=a!<>V�x��˽�I�_)�-��t���iz ����*����T�kǕa�Na�H��k~飦=/$Î@ 7쪮��yl��*�֡8��-��>����X?�尽]g����r�O.�F!��|��6̼��O����,>��j�=�4���@Y4(��(���o=��j"�%c�At�[6[m_s7�h�jF~��t��gTW��ηX�s<N�J	|�Z����ʘ�Ɂ�ֶ�"� ���9�&�H�=w*~�L��9�J�O&�r���y���2l^Ӈ�x�Ie@�*� A���;#�,5C��������ߗ�ecm�^��L(�
�W6�;4���aq7���lǛ����G(
�2|����[ѱ߻�~���ݰ�9zb݅*E�(����WM�a�`��":/�Ù��H��[r�G���[t=ز�)��3_Ő6���|�z��D>�������O��B;s���&�[(��h�1л�~�:����f4��4 ��m���W~U�b�����߭@��[�G�k��˝�T�nD>����9�93֗�A��*����=q��kQ��Gu����q�ldh�����e��/�,C��rG��Zb������:�����ȅA�!�4/yP+=.��'��q-�a��h�H䠟iT2��:��Uj�R��{PգJz�����V�.�!
�V�|����(Z\=����:�ט(�-@u?�f��|�%Cm�r�)���9k$8��\F<�C���/��?:�}Ls�'�}���K^E�����
n�,9�����P��*��P�rJ��Ѷ���d�$�7�7����4�������Y]�t��J� �F��B6�J�4w�U!��V�\���x��u�^�Z=q�":l:����\���.e�������gb�7�ݰ,��DJp��N�>4���`�E��O:G�үs�<gſON�2�1�5��5��d����f�m���}����L;m��U�>������0N�� {][g}�g���wX��1_���t:�r [��[GC2�E�*٨B�Y0P4�ɧ@�Y��1��_�2W�u��@��>�Ǹ3��<i:����E�'�*+��35Mp%܇KY�)w��h�w jB�Sw��Lk��M��=͝�p�ַ�4E{� ?�0b1�`���B�j
<벒G/�����3Io�<�h90sd��[L1nJPcA=yM�pFB����U�ǊQ�s �tj̃�� 'C�(� !��V3�-E� d��,?�f�g��������f��'�%.3њ���źe�e$z��o=o�7���M<�X<2@��,���o���E%2Z����6�u��]���4�0������0b��#���O��9-��eDu�������Tҽ�:�:âF��>2ag7��E?��M��� °ت~A��I����-�� �M����n������^�U
3<#���=e�YI����%�I[�Q�Ǘ`��HZ��؇$����2��-�����'��g$�{Gb�Yz1*���LN������u�ꔲ�}خ � ��l%>ݳ��F�ߨ�~܏BE���	���~�ө�)�V�W{��I�֟��+:���Py��V¡�L���ۯz� ss>+����n����Ή���	Da���bG�B�yf�YMk���n�o>�LH��]^@
��#����`����9Ì�/��dgS��-Htp�mQ���~i��){�9��/7;�� ���=��7�@θwI�i �fz�~ۆ�R31Ȼ!�UJA�b���v�`���ch$F����F�X�,�W�Sa�dX�
+z���!S>ԛd<>1��^��M�E���E�LR=��ʒ�H�ҫg�Y����
�3�h�5=��B �zSօ�;3�S̔1�LK8���7`�A�)��M��|C��A��-������!0��`��t��a��>I58a�������ٹ�t���a���f�����JGXY/x�9�03F��ӡԥ/�ڥ�9���|�<,�XP�҄�~K=o(��2�(D�	�e�7UU ���j
��7��^���םӔ~_S±X�<:� �HQQS�ۤ����;D�(o ��܃� SV�R�b�����}���E��1�s��n�"�C�i����)ͤo�,p�����gd�O_r�j��cڵ1&61T3�w� ���T��hu��k���.s�@&�.P9���N��g��f�.��,�b��ꜽ��䯄���_~D���tk�|��*�^+� +��2�(�z��_�JqJd?���F��b���!���Ͽz�|�.Š	�Ǣ�VG\�;��2�ՙ[v��5]}�����V�ߛ>?�����찥v���Q���3�w��`�VIS�(�S^�~�X�:a�~�������Lj����_�ɹ�5ӈ_[��A�����+�H-���7�;{�~���	��L出��Ε�+��|��<é+q����V�섆�Ȧr	�q(quT÷��E}��%!����v��'�C �I>����-�d��dXCM�Dύ�?�|�$������}X
�]9j^�AkV�I����FEn�D��d�vZT�m?��_t4��*�,~J��ѓ�����a�S�Bf���R���Ú����z9P��vʯ�Q>ƕ��ޚ\�ޝ��n�Y2U�?���f��,�^q�k�@3���>u�����eP�3�P�5{ߏ�512�%jl���9�;�Y
fQ >!<��1�Ƌf��?V�2�J9A�[��xei�H��+��mC6>l#���d�a��dͿu�\ �֨�HӐ�А�1˾l��1��O���h�VĈ�c�����ʄivC�A����(�Rb�uo�+�K+�^ꘫT/�������ǻ��W�;x����갃uט��&�g�룃�AS��>����;�Сg�SC՜��� 3��:4�^�b�@?�˽���e=�z���U�m�3�=�|�i�ǂ�j��cG���\6O����*���zͭ4:��̝%E�"A�����M�#$����˸��s~��@}\"�ҭ;
d�U$�UW��������Uud�7c.��j��
bt8���R�=Ǥ�t���7�^2����F��N�UΟ"[ C���"�N�����ߞ�8ԡ�?د?�{����T�\QZ�(c6j����.��n6Z$�����zI1�*@�V㇔��(����!�^-Q�W��Ǿ'_>ͺ�Fw �n���7�3t���߄�չk��4�Yww2�©�� 9��~�ɤ`b���n�S��!�,nf-�;4�Rf�f�� ��gB��@GGn#g\�G~��/ �	Yٛ_�?�����@=_���]����13�~Hxxr��ِ�0�����1�;w;C";��l���f\�#
��`�^D����.=
(���Kv�QՂC����g������D�(\�K-�{��am �RO���e��w��Wiđb_�ڝ	�W�wM~����l�}�L�-Fm(�t@3]zB���C���ˢ˘Iš H9�y���`�Td�O�q��y�#��)m�^ ����g7c	Cϕ�8�=�Y/������ٖ*����V��?*~v뗵�5B�8���yI������=�-��W�'��Z����z�Uz���J��( ϸzo�M)3�o��\���څ\���=�v���:r��k�H��K9��C˻ ���C����v���p�aO(q<�xT�UF��1�����͒4��N��BX�VZy�`]�2���S'�<@#���ι��Ь��w��@_C� �5�|&��壜����1(Vy�\�o���z���nk̜�D���d�mhݝ�+��=c�}�q&��E`��=���㛵��	w�-`��D1([܎u�x P�Meb�ؙ�-N�t2�-0?ڋ��!�۾�����2�4�'��hӛ���5�@�.23} ��s3)ĪF7��˸����B�QL�C-����@��g7�1q��z�_��d�.�B��?�P�s����}�Ͳqo��C��z�@w�a
�U<��m�6W�ns_9�s_�o�M��8�i�G<Z#U@�C���Jζ����7��kсX�jjp���a�Ŋ� QF����r4��z��Q����7Vq���{N׊ˡ��C����ߖ4�?%�����M��Fp�2�i���U����GbN�Ja�э��[����ݻ����x�+x!����T��a)e�5��A:jh�f[��í�Jb��;D6����������mN�6$*G��X��Q�Ţ��>��cm�o��}��n���К�ܔ7A��!��@��CV�5���E�R��/yG�R�C��!c�-\��pD�i��{rc���9;�sc(	;�&�"a\U��R�5cw�y�H�g��y�P��i v�60��I��OX�>s!�}����F�qst��a�����B�44K�DԒ��mh'+��\Px�l�i��M�6�Wg�K����-�������)s� �ћ�z:�!d�΍���/lF��mܯ�X���KO�D��ߟ�M	��TPY��g�h�/:���#��4�]~~﷡��>�Ϗ��ͳ�> ?�m��v�*�EVN��G7�f�ck�Q�������}z��[���*}��ڢ4}m��2����K�TF�K+�D��g)M��Ā($�FTa��~:�A�'���܋nCȋ/_�\�,��{��f_cV�)�l����% �Id}�%'#�D�}�����j���xԛ����t�̈́���-��RN��# p8�Q0���;W�|�����_��8�Ta�96a~��h4�L�(���
D)LO�<�tw��ڠ���ث��5V{����D��|y��g�b5PW�F�X�b��M�X�~�>�@�bФ.�{بЖd~�wĔp�C�Ib���y�lDW��y���7C�"���h��&�r�5�p�9.�1eJ�?��b٦��*���6�6�A=�n~����aqx�Ky�K�^g��u��4��#�`���J$W.4E�by��R�W�
6��Ƶ���"�5-���N�����4�m:M�Ca��ا�QS���R��M�]t�Oo����uGY�D�o'���f�Z��Y�(��/G�� J��Φ��R&��g�#�?���|��)���a�(d_�C2Ȓ���J=��M��r�c��^�Q�Tí�=�K��$Qzj1^?�>���V��� �3�?oa�Nzz�;���h��dY�!�q�U���!�E��p�Xqr�+\Vˬ����g�S�ݸB�����[��.�aAc��� ��S���������Vkbs�گ�h�5����G~�A��_r�08a]���!{cЬo���*�%�d��_YK��|�v�s�@
�����Kl��I}śW��J���|����Ņ@&%l��nǲ��A�V�(��=�pB:s�&(D�5ƽ.�����X���	ҋa!��FC��C_�1p��@�;{��w�e���x�� �?�8T*��=+�:�<�ka��n��Mf�u�u��)��
X�S���hb�I�0�<�[��g�b|�����Ě$��N��e����9�Ɲ"�.|X��4�2���_MS�B ޶��=�A{_�RC5�`�'p����������������R%�a^��<ێf��bre���
�a{��m{:B�m{�Ib!�o�@�@��R�G����E�h�j}�+2��NiFh��y�%V��߿�7�0��c�т��V���b�������}�n�"{`M`�rA�I�2�ߪ��9vytb����*8�g5ul��3>c=@��}p#��*h�J�9��Q^�K_������8�6����;��9�c�ܹ|g����웼����`'�P��E�.�/o(��WI���q���1�0���yl�/)�|;��S!�"8ֻD�9��Zê�̻Y�/��g6�m����I�n��0�>כܗ���	�2R�����4T�0�~/ƲX��%��nnF:���7&�O�Q�̡ ����?*h70Y�PE
��W�"z(j���jsH¥T"�SZ�k�����[ĺJU1FC�����o_*t%K\�l.��ݦ��i��VWHԫ�CU�����:G���o>�I�>竒�=�w-ג]��fC�|Ίu]��n�_����gt�I�n�"d��xt�7�B���m$>|��_ z@�XJ�Z�5u�趍����>���z�MQ$e0w7		�i)om~@S�=�LB7��X�]�<�� \�&�ң1�#��N0�a�c����Ӛ]��2L#��	��h��L��1�\�?>�cGEaGt7�����R���!6m(�y�T��y<��f� Ja�
8���k3R<��a=�]J�֧��d�_������ؓ�fYۄz�+=��'9�=7<�b���ɑf/l�4X��dP�4T_��D�4���*<�I������i<��ԟ�&@�H��3��|Z��'�� }��	x��M�/d�u9f;��� :������	d6s�P�Ǐ��e�E�f��Q�,�^������l���]�C���<m����'�����" 8w%�8۫��o>��	@ú����3A� x5���(�^(v;	�/$��K{�`s����I
�<��,H>�}m���\1�:��fl5�
=��9tQO(���^���Z24a�@'�%���#��E���#sK�oQ���NLր�Z�L���M(�T��lB��m�
����WI�e~C�c�(��&�.�k_|Ӊ7����򂨻������n����#��Hg\|=����OV2�]��c�n�)�`�s��n���f���}��`|�s
���lW�h�� =v
I��C�=L���&ⶌ+I��2��� � o��ӵ�a��Th�=i����?=,u��N8���e����%�%r~i�':bĩF��'����n��L5U"�$y��l�B�� r�,s7��9���Cp�}���Ai�.Ǔ��Q���%:�o��ʉ�s��˺�R �0O@�S�+�1��pFJ_��f>c�9�����\P%�/o3:�x�w�yW��&�Lce�#�	H�}w������W1xgI� ��|u8#�E�<t ���t5Y�kSЙ*BB��X�nQ=4�#��\�u�)f��VϬC��4�3�����l� �{��
�����Q����s��~6�<5�򺉗|���tH�;�4��jc�Os�
���g�	��(.1�Xa1���K�4���a�����\�͠�
 g1G�l	=h�H�� ��l�̖n�d1�{�X���X�$ٜ���� @�fT��
v����U�Q��)�W�׶�-y��;c��O#�s���m�Xפ#�*�\cH�
�4sW5>׋���w3`!�xء�K�����ǝ���aQm��艱^G��?���� �1v,Q(��̍V��5ޘ3��|W���9������l{i�q�%�������W{&�jz�-�An�՟��d����1ވ�g|��Y���"l���\?��T���JR��E̖/�3��7/N�`�<s�I���|T�ym���r�
V�Ć��c#>֍k9�S�S9#�����)׾��vۙ�r�g	���,�^�?����Ŧ���%�|�0����ckZ�( n�WD}�V�#P� ��d+��k�e��N�l��Kl��)^OH�K?]�ѭ%3�x��s�N�%F���ͥt�WsL��ъ�9#VB�s\f�����8|jt�ǅ�3���	D���Y��`F�T���D�N��m�7�C�`��L�ǖ�ޤC�M�}^b��OE0�"�Fj��5Z���Ռ�Y5m���!�%{+-G!��x����2<�]��6{}A�Hm��؛�oY�
+�?�٠F���ڟ޽��.{��-tʭ��I������z���E9����,�&X%�Ϻ*��-��7�L��pX��OC�/��w�:y�p�@��O���sܫ��:|�F8�4���/�M�i_��
�k�w^���&x���^�pl��i]>Ű@I6
^xn���TONL�MpJ��A.����>K��WSQ:�� xյ'�Xe�<� t4�����r+�	�7�G��I�C�B���g�mS��E���M�6F,~��e$�����	db�T@&b�l����["m��2m7��줞�5���	�4�Ŀ�O�IFDcK��7�rS�R)'�pOr��6uk��Ek�s<�`k�P�-�Y;���7ۜ��(���*b>�'�ڏ��'���<�zOԖ�N�l^��=�l�tp`h%���N�'�o�UH�7�j	K��9�=����ph�x_"c�A�&V���g@�AB��[�r�I0�c��"�2�I^ O${E6������r����2q���§�Xqd
,8�&KG�;uuy�-Ӳ?4�5��F�G�j��m6_-�K���]�
8kؕ������cT�lΐ-����"���;��BY$�/�-ｰb�i`���r������FE�:�-�9*�>���^FK�5���i'2�/��S����ߣ,�DѨ�;m�cs$Q��އ�o[��Ꟶ��%�*tS`�--���%N	1ڐC��|��������Uf�ݽը���{����f�Wf���_�%��u�7#b�����xc�4��>@J���-��Y����@��q;Z�� $.�v�YO#�`�v��(Z��1����%��0��v���ks�'2�}��e!���$iB���zN��6��8t*��
�Xush5����y�7�r�
  �˕���c���L�P��(ע�����3�-f`9��'o�.&���0ˋC@����������U�b[5���\�G4���ՙ(�I���{���S�#���t):ٝ��)˛ƍ���J}��WYMr�uC_=�0Bv����ݼ�����H�P��_��">�d�L�Lr�Z>���	���#�f���*��V�?kP�{�l�zε�t��%�xi��oeȶw��O`aG_i�)G�$53;���|���!�����.{>����2̈́��с�跎�u��L��שu�kƻ�K���u�Ё�X|B�f��&oZ�-x6��l��5��F�;LKi'���M��߯ܭ�ח����[6�#�7�2�Ikb�A�D~ڈ���}'����l��d����ie=x��-�_�K��Y������LK2��bb�s�*<���v��+��c��<qj��J����]��5�hӴ7{
��@$�{�1s��)ۃ�&*5J68ql��`���Et�f%b)Lg�ۥ�>�� �e�jb��Z�����Mu��L����pl�M����ٗ�)��֔�ǿ������C������_*_�s�k����rO�"uq�7�E�g���%AಉvHF�d�*��$bq}`V��@l�$�j������-�0��a.d}.���I�ީ�Q����C�_��5{���2|?4;��j��UQ��i}6����R�@���+l�{$��.��|��#�:�(���q2��Tb�ϖ�ͶWe���i��`<�>X+�Qe�C��ȣ7�`z��E�|��|s�/;d�k���5`�ŷ��0��gPE�V�k�o�3Ǻ��{L`e��S&�ϸ�U�d�dp����L���(����cŏ8��ʎ(c+�>$�l��7�7����������x^v�p�(�!��3������ W%��j�F�-;�P�ά���3*?y?���jkYs���I�sե�=�R��h��A�[��Z9A��D�1y皰1�]L�Ts/��4��0�4�"̷^��&R4@�	
��VD|�p��E̋���q�Y�'Qݺ�X�-��T%>àA����%� '����ϣ�j�&���ˊ�.�x�>!�7`� r�C�X�O�eʑM��o�5S�h���FF�-4�&�@�k7�Ԑ�#���� %�R`\Pp���z��\��W/6V�4U�Ƨ�U��+��b1L�_���  [6EgL���@������{Q��¯�ȍ�O�6<�R=P�ף�{ �r0��B��q P'��o�˦�B���W�M�!:�K��j'���ހ�`,��(a�=�����, ���âG����:�"��>;[0�7���$�3���T+���^�#"� r�ޔ�1u��1��U�p���%�9��m�yL+B+��uvu��.���&
�J���5�{d�:���O
�i�Bm�%x��I{�F����U"H���.}����ILד?�R�b	\2����OѣK��&ل�����j�e�"t켶^��4�vF���dbT �+>L��	m�) ����.&�����x�5FUߌQ��n%��%�"���������ku�K��w��5�`C�&¤z�:[+����}q�4��2'�
_����'
7��H3������Г�޻��p󏯐0H�����Q��ܞW�v��1���(o�h���d�Q��.��__j��}&�J�n}ٛ4�sL��]�����?��UU`���)��R�CF��D�n��hq���f�p��z�Q�4���9�Tn�A��}��h�,��g��j���:�{�?��Z#��*��ϳsV�&�aT��f'�9��%5� ��nhr���G�C�;.F��J�@iW���0a�`M�y?a��Nar��>ڇ�չ���X�$�H�V�N�Ѳ`�k��-�[h�:�8�(r��W�-��ڑ�C@�U���o|�*<���6�"Le@�����ݘ�eng�:8���;��	`�P=���/s}�/��.���H5�.~��%�1�ы�'Vi%�M4o�"ytјe��)����c�ޢ;���AEl&^�Z��i@Rʋ�ܘ�_���S!�s�.W��6�)4]�4'p Oyx릃[��?�1���@�b���:��� ���5�d�������ϔ��F< E�VnL"�9h��;㎭�{�pt�����]�&��뽰\z��C�b�J���&�8z�o��y�9�w(۝�Ԅw�������IU%���Ҋ��fx���w��{f���^N֎"�tCUӜC���$��TjAk9*��vH��d��z�;Ң>�Ǖk�j������F 0��l�����	�	1�B�o�r��8̺����B�t��4|U���� ^�(�U�5��u;�KfN��(�Y��J����*�)���[�-{3�hU!��S�[!ؓ5!��?�dA 7��/��%�Ҋ&�͏zK����/-�Wd�$�Iն҂�����R����(:���C�Ğs����Y�Ԩ,��/=$�S������=�Jߣ��`~���]��J]��9���\Hcf�Y
,cۈ�|����I�)ySy���$2�-�'���n��[V��&@+,W,-�8]\C'�~�rO�ɞ���S�ǖ1.m6;�����{�13��:�=�'�Ӳwd��WRF�Y�i�"w(e��� �d��ǫș�ԭ�
� [�q|ɑe��{��;11>�_I���������<#�{��q���mgdƅՠ���=�v�y���f�`��.�W��ɤ��{��pZ=���%L��~�2}xe/Gf��4Vi���q�m��i7�6W>�nN�w0#���=y�e��'5D�-F�7Ŧ�A|�P{�aX9#?�Ch�M\���r��͟��W�Ays�������p�& F�������a���F���ߦ{��3�W��8�_�R�ᓢO���Va��ǲ:�T��"��¼L�^���7�ΐ"kfGO�ӧWa���R�V��S%\��h���{J�y 4_m��<->�né��6���"yHZT��w�c@���m2�.2�Hw�$~l)p��L�P��Uɨ���cg���gZ�d��1��a�X�^w:?��sz��uYE8�O�в��n�o��(�:����DO��.���� �u�Q�}27.��4���9����"t`���>��P�H�0O|j�E��5������8����Z��u�ᡓK�@,�4��_��M�{/'�7Ԃ��v����.�Lp����m��p����w���6��X�[[�)�E��\i(C��,��x�oI� AM��m�p�L�嫚>\�y�T���f��1	E01����˞m�/�PށF*��B,-�/��ebD�����n���K��r Ud,T�by�r�2,���&���%Xm+�(%���m��r��4�e��Z���QuH~�&����s�����ѥnk�=e	��S�%��k$i��S��d���$g��2> V�-����_6|�\��;U��꾍���f����^�o_0̋����w�H��yP����ʮ~ބ3���;,}�Ɋq��-���.Щ[��?ΟPaV�fd���X�"γ,.������ )��u�I��Z�(�[?:��P��b�Z
O�a�޷.�l7x�H��kS/�����G-�`�C�|�_�W_�H��f��I�iD�'#?H��yb���)K�/��Y��mӏ�j�Ͷܤ	���-��w�s���c|z%�1KnK�Ӣ�Y'v��7�*l�����62J�\*T\Fr� �ir��wk��@�E������zD��F��D�<�!o�*00"�}1��z��8��P|2qY�\V��z�d�wo�ݷv������_S���ǐ�m���.�q��w�o7�هt����ЕS�S����d��BS}q�I������0۷55ɩ��M#/�$�@�`t��I�>�T���v6��S���([�
yNP)b�*z�Y��J���G�D1�|�g(��� �#��mgy��a;@D��I)��ZEa���^fiaf_X|>������)d�%[JB����K]/9�WEt���,�J(�7�j(���i�kT���qO'D�4�XX���:;�:9`������o1�\���C6��S]]�����U|"
y��ZО���LX�'�G��`
�a�q)|�t6��X0�3H�>5&`�p?���y�LJX��L�\UG��+��1Q�3�x0b\�W7���a�m�@M ;���#3�̆�vcwR&t�1	���V����Ud� �� ���U'�dhhbD 4�/�`��΁F%����bI�պuB@�&�%u�Г�t./` :�wY��Jg����ef�D95d_����j�\��0�i�o)���h�	f��jt�)�"r�o�����q���_�#]������/.���7&/=m��Ut��/+0�ϓ����~���.�����<�	̦x�����!M����zR�s����,���N��]��Ct�ˡ3Gf�G��3�q�2�ri�b��rY��5֬y�4�Gk޴z�^{ ��ry�����a�	Jg�f4<y1����_
[��(��\��`�f��ŭ]��&��M�4�=þ�AV���\[�]�n>�}$��/���(��mX{mG�ˠr������:���cT�x�=N�#(�E�J�BX��b��쫲����� Y�X�]g0ҡ
J��{�{	���uݞ�ʛ�;ۺ=�r���X��ꊕRcH�C����^��O�I�q%� �P֐�*�D9Q�jL�U	qI��`D�?�>��x�ժ ���L��3�Q�Ͻ]{�\��Kb0�C�5�'R�e�ܸ��ڵ��5 ~�y#�Ē�q�x9�#YU阗�:�Ν�,�y�j�'�x_5���cjʘbR����At���Dfl n���0o(��T��t�v,����pm�B�%��m����&Y7�e��f`y=��gn@Š��<�����iU�	�Kb�%����a-Y��\A�bx}�r{#��w�4�r�.��! �Vvu����1�n�U̖x�� J)�$�!�֕�,VO��e�g�š*�^��w!���>}�G���������q=[�E�m����pR(\��U�uv/8��M\I3��������n��&��r�dq���縩dpX��s'�e�5�!�l����	�/.)�*��8Jo{ ���ØW���C{�mq�hy�:�Y�`�b�k�9ֱЏ-[X)_~�����Һ;�15��d��1�s��[�:���g��7���u�{	�A���o�a�uo�x�MƢ[���ټ���99��u�L`��� 	x��`qIy�ƃ�ą����#[9����� �tq1R��"v[�n�R��-����d�e0������ m_`�`��(yq�$jH��Z��d˗�4r��25	!(�H�� Y/.-���>��}D�Ja\=�15Q��E���y�M�b/��b�ޛ���y���ĺ��� Mi�`/�z�/ y3��ř���/eѲ7H��r)�8�S �}����`�9P�Ey���/���D�	]�v5�͝X��I�X��]-�+e��1�8.�u9�:��F:��g1A�lv��M`��a���X�� :�~�u3�.���M<�7���^��!!`c�́���2�1w}�8�) �zU=�B܆�R����m#h&�/�3,v�r�Z51�(,7b�L���O�?�sg%�leW-�F;�|B�x��F� |e]�ܱ�ǈ��6�]�sʮޅ�� ʢ�A@�7��+v>E0_ZT}p�/K2��k��1\x�.���|�ިv$�d�GA�<5��K�=JJ�Vڤ���{��x�l�B;�_`Vg����<Z���I��1�#ͰU@���J���e��C[�����	�M"�g�� J��+����B&U�LOPQ"3���xz0Ԗ!�����v�С9|���w{x�<.���'!�$�(5Gd��U83�₅�6=JW��#2T�ʆ�h�%6��p�#�����0��n�jm6JS�T�	VJ���<k����ݞM���ע
{�9��y��Ύg�l��((_Xx�>CY�����w��:w��x��M�@�������sy�N��Qja��r�;~M+<%}�1x$�qY]#���Ȣ�G��K�jha�|��%���$�|��8��ߎs�5�����Wnš"���6.���(y4���{���z���H��̬j%���]����V!�ղՓ��5-t�����c���G��1���|�*1:'���Հ�>�v��nAa~WO�Or�����ȹ/@/X��_U����ْ��qu�&B����˓ftժM$a\>j0ɼ6`��n���sG!�(�v�I�c��YW������+ަ�tmӆ%�GRA@\p������+g��hl�����|�t��l��Z#6�R���C��鄇� )O��@�~����I1��d���#���/�����٧�2b��1��%_�5B��-��5Ǥ����<����중a�"v�lQ-�g�;��0Y�y�c"'�CE�����<�}�G�? $=tW��ҋ�<T�p��yN/k&ˏZP��41Z$�7����H����&�k�>k���N�]sI�O�SY��f����7Ά���U�k���@�TfvD�h���7�L_C%R��Ș�YQ�pH�=�Xؐ����.��a�����M@�|[�eU%�E���ʩxf��׋�[LDy��y�IH$h`����'�����@���]�e�j�m�}�t�B2�"|�/_���M!���(4��l���3U�B]L��{Qmq���rTT���)}Ջ˵��_���]��ɍ�i�i:����vͰ>��eR�m�,�eA�U��K:�r�w��@�̹<T�Cw��	.����gEy˱���J��^�ƛ����˙�m	���*�O.�"�y6��~3�~�y�'�K�l�hz�{��y��ܤ�&��R���V�2g6&����Z���[Ƿ��[�q���5k�҂6��R�b������F�2�>�ĭP�ѵ��*Ƽ�xQj�B���g�M��b��[JpԴ�=�#0yp3|�X� �_�6|��s�����%��o+�����B�Q��Jj#�
�lZ.�I��HE(�z�W΅���B���O�]��Ȱ��	A���P8����f����#Ox��ඌ��畾V9H4�����u��(�h)�05C)k!�M�6o#2s�nW?Kj띸 h|s����(	���H�*�W�7��g�K�c��xV��ho����w���~�;�8��x�0��H-\!*�Ԧ$�7�$�^�S�|zF�Yߙ�n��?i���,b|-P��5)�M�ӡ�T��%���C���
��M1�YkJ��=��03���r`�����x���wh�_6U���˭��ZC��呺:��������)oΑ �5���v���s"l�Vk���r�qv��t��H3iW˃�\��wRSЃbQAW�[�&�0�`K�z�w35����EYWڥ�fq�8���Ut�>�(*m �l�D���w��)�
����r�脖�L�g��l���T�	��a�����_�WU	c���\�h�KE4tz/� �|���f���;:�%;�����9�q |�8[�z���Ӱ1��VJ���3���r�A��w� ��iT@ 
����q��ƛ�3�-�����~�ׄ���Υ�megq��{�@h�&#޵�;J��H��7�S]�����굽N����I+K �F{�����C�����A^�GS=��2W�j�G�t����je�U
է��jl
tS��uY_��3B�S~7���E�C��ܪ�fq�`&���C�� �'��A��j@�� �/�`�JQ����H��0	���)PM�#��aA� �����P��,&�TD/�Wu��"���������()+�m�ν�H�ԋ�x���a���J�8E/��������9�;�U�0���3?iL1�#��)˦{�YOn��sJ�<��Nr�ӕ���	X4m:K-Io�yMJ�쪨��=��͌ԇ���l���Eo�k_o�w���N6�[P����4�]ytƓf�iBa�e�@�Yٷ<K���a�P��\�o7���r|3�P9v&��`H��s�ֻIj��L�f�h ֬~����?L�^�K#�TW^J�P�D'�PL�T�"�g-�r1�pj��H� �S������E��w�L���U�����(����tɇ�&��;�e�A�+b��o�^���0J@��ݜ�����5
^�"jh��Ȑ�A�x>K�F)���ϡ�D�:���}vT��1��IΆZ�)���#9@řg�%pZ���{�A����ڠ˥�T&B`�h�És�#�=�5Rf�����|o���
�����/��`��C$�K	c���O�q����c�VrA�Ǽ�b�b�s��)q��狤���H-'�7w��u�	p߽�X�G��" �9�>KZgH�9���)�Z+�|>���2�|���ZŜ�&�P��eF)�ú�t� ;��h!�M�x
��p���<�A~��Ir�Q�Z��x�N���������V��x͝��:R��ܮϪ6��0볎�F�P���A�"����-���nM��E<a�&��J��h��w(�.M���
��÷9{���5o`�����X$�� �"aH�A�%����08W3%�^4��L@���_$GV�^W�#Tw��W,p�V6A̴�J.XQ����FT��H�?�y�dn�s��ct�_ýȚ�:*"�qO%K%�7O>!w����y ]w���UuҌO�P�΀�,�ɫ1�=��]İ�vBy�KJ �E-Bf{Ia%�c˫�����ٖ��
~$��X�>��f&L��5��
L�R��B�!D)T���"��a��l��Du��f6���{Xh�Vr<�����8�f��/Ͽ��e���3�_u�Ưd�}���s�tK��;OFP�/�ɮ'�Fh���ﯦ˪h|��)�@0;{�������+�F�+�<�A88w2�	󛭽�!
�3嚺oV��&���hC�m���}��nV�D���kEv��{�k,��/5�}�U��OG��7�_}���1���YL�4.�eE���脷�0+O
ʜ'Z����i�^��b�Y-c�8\l _�g[�q.�n���MҨz����f�NR�g��\��ݎZ��^&��S��*\�9Q鉦�ː�a+�2v��.��T��}���a��Z����X�k87��[.�Jm�K�i�:X���5U^9��p�ky��L�fͼ,W�7�WH�a����ؐy�"|�=����z�ı��^���)FU15�
�=�3:!��D��`�ܒ�܋0�x3l��QNZH^�8���:cH�f� �X�F)x�ё�4���(��:��o#�:kf5�����Ix_"��;l���)r�X;Jr[o�t��qk�nPB�!W�-<軃��94��A�2/3�ٙ'���`�ʉz��ɝ�E�n�%"�*sLiq�V]?��C_8���S���#e�;��ҝ�jI;d�k��\�Q�>��2�UX���*�x�u�AA�1�HnQ�U}���M0���Z�9��p��'��oQ�ռW��x����K^4N��� 5GV���/��B>���Gr+R�����Hr�@QN�j��u$�؂�:��u��[�YWE�*w@��j����̭*ؚc���9^+t�E(Zh7�<�Ƌv��T]uN;����Wmwx��]*Ʈ�==<�ܯn(n#���VȞ��'�n3���M��&v�&���h��c�c�DR�_�����C��7�1<�1\��T�J�?�S�	T �6��O\��r����ހˣ`ۆܾp\hﶘ����i�Τ�ї�A׎��q�Y�A-���)��:����R�u��2u������-���=?燏)|�p?湙�u�w�8�(�գ ��7�N��*rv���5�i�:��)��XZa�3���o�A��>�N��t���?	�:��}&"�Ėn՗[ص$�&�j~���}cY�8���J���wlr�a����Űl�S/z��g�\�x>�FIse�u�H���!N	s`�U�����b�*:��0�i����ӑr���,,���eĢ�F�z��QWN$�S�����f���/��'����x�޲��2�ҿ4��#!����Ɋz���O��_(�W��kT�n8��BM*|�F���E�)x\���n-�7 ��U�L��h���v/�D�����ϡ�����F=hȾ5�p�퀸�5�ՙ�IJi�L�l����x1�K#�6�M�ǟ���t�S,�ŷ�i_�ZO������>.�P��G�i�R�.ba�7}o9��%����oG�_� ��%�3jx�j+���3e����-?�?3��l+�6��K8.ע�=�v2���~��iJ=����=EE2y���#�&LZCm(��h���}��S\�Cf��R�#�0}���B��KER6^j��i�����x�۟�cY������Юy����s��+�� ���� ��"b?�`��w��k�n��z.m�ed�7O	#��i�T\޶��I؝EX'��������9�L�=��2Wl6S�K�_��0��WJv)2@(D�*6��O���j/�c�-�el3啶jT��[��aײַ5����-=��v�1���C�l��������(d�S*T�N:�,2�I�KW��1f�M7_8��m.���U�ZR,w��L�"��[J6�*>)���Ybl;����H+^�YA��|iI�y�Rى�V{U-�4��#D�B�k�Tw��LZ�"~i�@�3��g�nNE��p�n��u_[I�;%�3�Vb��@��]��9Nq������t2��4�<j �X�R��U�s��*
y��!߹RA�C�����ݘAeT�A-y�B�%^�+��9�)O���
+7�n�ł���2ֿ;ÔT�=��.,� ^��<��O�\�[�� �
��D�k�P9 ���c
R�a)1e	�1˧�&�J/Q'X��3 d�"4�S�����.R���u7��]��7yD�^�&��D��C��̧�S��8�Ezn�MD���	opK�BQ��7�;YO��R�^���apeN�l����Y͟���Be�74�^C���F�2��bYo�m=���:q0K?Z߰�}E�1���pe(�7w"���gi]}���bW\�$�]�7�X�L+`��MI�]����;���S0��ͦ�]����@W$
����I�0�O[�����P%=z����&��ϛH��>Ux%E�^���ɾ};άfpY�,7:]d��cA����1Cm�}����_����@���C���J����"[���ӹ��@�D�	��r����E���Ѧ�'���d�#\�=Q�w6��N�I�1\��R��E�f�ܾ=]�ؖM���,�ύ�f��+SDh���_�@����9�H?J��;^���G�������4����L�,�����з��:�Mϛ��%���;2T���Kzsg�:��I}�ɼ��_Zײ4���W�@�cN	\�u-��-a�}J�Yu�����)��(H��Zʯ9v,����JDʪ�������t]1s�<r;p�t�N5`J�2��ɫ��z�cm���%���M� �������z�0���暅�3,-��\��,� �*�Q��	q�����N�sJZ��}�{��Wi�\uF��g�'���̈����P���R���m�\��b"�D^6�?�>,Vz�&l�z���|�l��V���xYi�D�KSM;6���Ĺ��aa���)8s	�ޘsC���oi�hM�c�׹�3�~�G1ފ����4���l� 
�D�7�9��t�xkO�ٽ�4�<̟=oG߂rv��a�;(�p����k�)�Q��kz�ul���{�lVӔU�\$YvC�J\۾�����0�w?�v��Rտ�D�����w������77��](o�F7L�0K- tl8��׆�d^���'�w�s�~*X+���a�7U��~����ӼՕY�Ѳ�$u�_�fK��F��W��9����X"�д�u��Om�9�P�J�q+HYڇ>J�8���0ˁ�v4�"*>��������!0y<A���\�̀F�9!$�:�e��d��׊C<�t]��,q�1x ���(CA�l�m��,�R�8�b��`�|Y��a�a�����O��"�[iSÄD�V���H&�J��6�ܱ�5$@�o�"��Pr������rc�B�G(r�r��;}ܑ4�(_놃�a���!z�ש$`�I�+��u-L�@(�q��h~T"uɶ���C,"ssk����<�7��^|��hS���&�*�A�P��=�}���@o�kw�<�o훀��b�������x�º3��G!� 2���(��;���E�0�v��Q�|��G'�*����&��
XG�{�08�����w���Æ��A��pͦ+m�A\]��]_��Z7�X����:��.j�M��3j�$EN��n]x�j��-C����֘7n�B������㯵�	EN������ a�dK���G �v��L"3�c���"�`�:�BqQN��?�����>��H�JXF�4�y���y��i��`0u�Z��O!���H�4Ʉ���jDc���p� GS%��"�e�M��+%bO6T�u�TX��A2�,�u(;���L8���_ʆ?��c���T��7����O	��.vE?�f.Z��t_�z�Q*��:o�_�j�N�+]	�CZ|�Vq�	��o��&4 m1�,a��X ��6�'L����1
˩ �,H�K2J�%t���_k�7q�*�M���2�!h��f�w�k�`��AZ�9����R���3�GJ��Nm��Zp$i[�>�������/��^���h���,�����p���.�ɥp�˔�-��wo�w5��3�/]÷��ƯEM'(���+�C�����ju���WW��1�W��(�0��H����0Ն>�(�oC�J|&=���%\��U�y-�e$d�ZkV��r��0���U	���O�]�@/If���#����;�F��ԯ��;/�ݬ�E�QVH��0R�$���$Q)I�g�\�+ p�.��޸��cB����L��z��/�J;���I�@橍�6�U��e	Vi3˕=��E�,�9��tU!� O���_ojB�t-{$�5L����� �gC�ѹ�ؽ.u�0
�CK�-�6^VY��yM5�~��~�qhع���]�����U�*�A�N���a�,~`P���M
rQ8랟�����bKyNk�B����!��ϼ��P*���A�Ǳk�T��zQdeҲ��|й��K�q��3H=���X!���:Z%L�Q>
�}݌/�#S�9i6D�O �KP�nu=W����%�6�����z�=��j�qYm�t'ß�����ӕ[<� ��a�~ ����&_=�T���X�W��x�w��5�����a)�@�=�d�h���a��_
�#E}L�{�������,�f���岢j�����5��a��ԉ���l��7=�r�yv�t��%/��8�v�0`����	��lRA�7Q�v��� �^Ȕ)�0g�f��y��fw�uL?T���sq�� ��w��e�\`\E��|?B>k`�A^�#^�`�(U����[l;<_9p
�&����奫g���I ��܄� �Pb�c������Lk����Ǧ���w��!U(9h0,��Z!�iU�l5GJ᭯mF�����5��w����Kir�{.���O����T?D(��H��S���N�q�l��};*����&dVp;Μ��j+U�ɪŪݧ�2��|I�4�����쭨g�}8�M���xF�Ol�k#?��?�Mo�D��o��N)s�$*�e��SgTt+c��@�?Lc-��p�Y��B�hC��o�[�B��]�1�x�"1[���5]U
�".o��t-s
�k�uy�Lt��D�7�jS.��̬Fv�դ���ʺ�����C�)�Q�V �����Й���38���� ��,L�E������4���A�V*sW����ޅ�sZ�y8 K��H�9ّ��_�	1�pg�u�;O���e�[�bb��d���2"Ü7G�Q ���q����ˣ�:}!���@|!�&�r�e��(b�f�6�ߙ�\�rYd�*�ԝ�eyQ�f8���ȋ�w�$�O�������1�W�W��FB�D9�����Q�:\�=R��1����N�W�@�vK��`�!I�F�;Ί�:~n�
n����0�@ȥ	x|ѱC�_�d�v��O˯�{��$�^<�yAhڧk"1���tXZw�:Yv�W�
�V��}_��'m�k�y��0�1���EBea��Y�$�eh����lu*��=%R
s��C-������bg����U=��R��'�7��#�Dy?��X���Q�$wX�4o4`mM����:���U��N��`ק��u6m��E�J
��g�c �=�+���O� |^������>y���b���;�F�P��L��TĊA��C��m3a��$*�,�a8�q���-��ڮc}c	@�<�����w�������z��z�)bz���D�� ���k|J�\>�|��K���C���нe+]p@-��N�<k��)ⷽӛ~KN2�re��ʲΈ?��s�!�p�I��PE���D�s���x�-	�*Th/�;˥��4I��U��"OuCA�oyi��b-]����R��B�c��v=D�Z�V�Q���>���΍ln,��ֵ!��cE�����nz�m���դS�*�R:�A%ʿ�3}5/GxB��nP�֤���k��&^3�A`�v���k:"�o�����Z�^���⌣��~��1b�ѲI�3]3>$f$<����T�^�To���=���fr�H���_�l�M^�ɲ4p�k�ؓ���EX���_ �d��ٴM4J):��@�i�ݲc.�9��?�	��z�#v�w��&mI�U����L�N�ʣ�cj�6"Ak=�=+o|�Yl�x�*��RIVO},�@6����1�4V�E�J�����K��-h�<9 \ST�8��}������VՄ�G�u�6lE߬����$�X�U$�E�Ț)���(i�e�Ʊ��-Q���{���DU����Z��<����$��gC�p<R�N�a[������m����d�<%���M`K+t�L���_���Ϲ���,k���$�r�i�W�v�c+�0�/�᠈-�Ju����6����d�Lj�>�%�YU5����^�e��3nJ�l�����c�z�Ț�p������si�]�}/I
�|g��B��B���5u#���J`��+D�_�V�t�X�޾���e���++(��N���7����4hF��Y�`TF(��[B٨�ܲ����j孹�z$E>�1�� �Pj2��-/!#'��\��s>O����
��[�)"'M���)�{��j!�Ylɗ �De҅�~�$i�ߔ0b��M��hDv��2��*;��u�y� x-a��yF�����^�����m�㐉Ԉ�!���g�\�>+C/{�[O�k���7�g�Gs-m���Yi�g:և�b�L�h�q��Fi�3�D�����OJ0Tj����%�/-��I��Jc��W��C ��s���/l^S`A�~h���"v �c��DE4�qY{P*+c�sM���L��J|���6��f0�40�G�RW��G���R�&�hB:���ɡ��;˼n���֋�,�m��}#~�+W���챗ĝà�<S�ڹ��������L�|���>7����w���i�@�15p�	�����u��g��3�ݛHY�m�y�x�f�B�e͟#�6/Uja䄷/I /�!_�FA1�)�B�!h��eW%QD+dZ8�A�(���re�[p���<��ΨN�E8�BD'�vXQY�6�x3|��V�F-��s��Id~��:.2f�K�+%����������M�?a�g1���@�a���	�D��)�R6˖\�l�(CN��:m�j=R�A��.�}ڠ __��[�Ř�wb��}��Z(+���gi��&rQ�9����"+C�?t�\���(���f!y0��n�S��9���B�sl�@��CC�����ȓkO�K5^�%ں���z�gJQ��t��T�"f����ʥe3�J���o�z�QydwF6�n��&�k̰]����^�
)�6���$S�ہP56cV`�?��_�O����MǛ9�d�"��b<��$r�3u��wZ&�&*�B���x#�uqۤw�p�R2��;����fdFIº��
�҃E�Ɵ�y�@�#tψb��K����¸̎�헿��=.W� /VX�L[�.����gd�jYA*���,�mA+7nRy�KjL�|;6<���2c�MƗd{��[��TC�E��y�w���ʱ/�0C�1��:�ޱ�qB-���w���
(q�nHQ�=2l l��}�<�"˩n<K�E6����h��J4]E��8j�FB�'iZ�3<u�i��y�G�N���+���6����b�vͣ�Z��ˌ�d�=��N.�"�'�Ju/�}�R�eVe���)6~���	.�'^�X�f�AY��8Z����B���eO���1���ԏ���Gϸg/Q�{���(/�0W'<~u�L�H�u8ض��7XM���6��@$�-�O�r�i"�U����p�R�����Δ�E�'^���\��
�����g�P���<Z���ڌ-�<�q�E%�}��G�#��iۜ��A�������Vc%�t�oS���{~��k�Pw��Ƣ�d�>L�'�і�Ѕ������C1^�w\S��<#*�I��(;Jc�=Lޥ�X:��i=@���*�Ւ��D!(ݪ�133�9��a�w�X���
�׮�i4K�lR�s���ٻ�������ڹE�$�c_ U��+/�a��4�!N��0G�J��ܬ�I���f���)76��L������iʹ�Qx�I�d] <p&�x�n�D�d}T!d���<��X��p!<@y��H�B���`���[��69� c��-��\7�'p2=g��>�n̙��ECN�%\�$v�_@&�v�$�|���Kw���2g5J_/����CF�Vn�E����^�ď�ڧ�/W:���;�hy3[�^e�� ��D��ؑ���z�q�Si����{�䗨o����!�.a����Z��͏cca����~8�
�pY=�xR�!싉3V㻙�1���+<��A��
DOLǥ�U���ꄡ��˳�GŽ��&���j��(p/��O6��:��n��Y�����=(`6El� }���!�A�̨|�E�5�a$�(�0�F[��5�k�u蛂�
H�W���C���
����K��2�y�	��rջ5���MJݔ\zʬ���`9�~x6��
[+�f��{R�� ��9n<F+%�	!MrvH&�L[�uB;��N3�鳿$�~�x�p䘙���JT�<��̖ͳ��½����9�*\��N6/p�7�ڮ�7;�r9$~ _��f4
�#���w�
%��Hv����a��� 	��ܧu�?��"2���1vhz��l�
�&��](��|K�����2,�s[W+�@� 6&�Ct�7�[�k@#Wd������3EB]
Au�ET���q�[�6�dbSx�:Svr.���mg����s����t�u7�����w��*��iR��y�ZC����?'�X,p720���4-j�lk5}����y
m��n�m=x�J�\�۝�M�{�N-�8K�ɤ"Lͳ��[]���r�W�y2�4���~*��ټ��%a�7`L>��*������g����\F��k�v�þ�d���Wn9����؋���i�0�C�	hg	� j;W��ù뇒��������X��5���`� '0&%=!�EP}�+�N��n����]P�S8�ĵ.opH�cod�8||̹���A�NV!�?�Z�B�kg��l68�z������H,��O����tC9t][�:P�c&�e���S����H�������)�{%A�_��M�����M���&>���qA�%]�mM���t9��t��(7�וϱ�Ӻe��FU�@��\���䥽�1r���@.�]|����Gs��NgD����ߊ�������T�Ώ�#��x�٬?M�����q�ʳ��� i^ Ơ�˙M��	��Ov�4��(�y���7�1ւ�x�h0?�c+�_�ZuA"q|�
�����o�Q��utٳ]ŦW��+U��
2c����T\��5�Z4�4�2��G`w�������}S�!��R�!7:h��-Zc��H���h8�Z>k��ra?�H�ߣ�C�BBO�,o
�����
�d���w�ѢU�
-���l�|m��,�Xl=3�Y�+I���)E�?m�ӝ:�y��z�����k�����������}H�0�~��ɃqM�m��:�+;�(n��&��q��ƾ(��W�qBd8�d�{�4H��'$��ߐ�j0�����כ����[K1"G8��QX��L��fs��C����}5��_��h�^"�r ~5za����3��1���|^��u��р[�(��c4M����}���c���_f:������8kl�e�I�zn
-�MJ�����m2xm��'�b��]�4��!@.�V�o�j����},�TŧM��%�H*�]*�����@�k�2)I���j�2m���J�r��A�?�l{�����/�v���C�_��Ux7�&o�n5�����&Q߭�"��L��=�L���mB?"�J�q�������!W�2Z�a��b�[9H���jߌƹVg1��Ӓ�����v�3h�f�<|�&��`�0���%vL���O�%A��G02M���-մZ9�Y�������B�Q(g"fo�a!q+'iO�w)/����T�s�6b�4��������\AZ��2�X\
M�%\��	[���Vq�]�~;!������&>�'�HQ������8r� �*�z���[�g9��$�"���c�=���w� �����?�g�΅���RV�t�� ��K�h�ߢ�Mͯ����Æg��!r��>nP��u����/V�J[��lw�	��9<�-Ry��y��^G�����h�/)���z�؋@������{j�pK��66�����6`J��uX�:s�=��l)�]�IV�۠��9e�p�^F*;w3��
;�����N�Qy$��Y���E��hG��R.�/�i]�[WV�o���ja��nP?���D�r���۷�/�<0q*�t!�;������-;�z�9:DB{���x����Ԉ��`��4���8mm�D3
�В"G`�tؤ���lK�̎t��W��Ŋ��]3���;��TJ6C!t�/Ks����l��$Po�~���������2�]��MU�6O��4v(j�T�X��JPRB�:)R�݅Q�~`r�����
M��<�9Il��mJK�4R7)�������f0QM[h��>��&5k_.������@�54�0���̒�s��F/�2f�P��d���A'K�S�L�mY{�*=�'��E�� gU;�����>���|7���NU�p�:������Nb#ZU�f�jC�u�ӿ��c��kmw�wL �4dJȓ��Q���Qc����z�T�M��DL}Jm�k���I���p�6���=ȵf���{\ dBh:�>��佰̃�;��I������{��kae�+\V7LZ>+�aϩ ,�w48�I�P�c�4ΰ3v�ٸ`Q�_�H�H���<��L�e:��qX?�G��  ��p1#<�ܻJ�&�$��W�g.�����5@�BGm��F* �ÄhNE'<v�����WZoUGxƩ��u� r@���D�x�? ���;y�@�Ie� 
/9'��QG ������=%�hgf��X��(J�ԷEսT�nJ1)��oP:��so��@,��9hR>̬R��;��9�۟j�?�ai:�S���$rZ�󄣡F��<\>�~v M�Αi��>�-mK I|tx�bڳk����U�H�Ya[*àk���Mgy n�nYlf�߯ଁYS�*���Tİ#B�u>��(Bp��5�C8��4i�܃�� �Vb�П�81Bw��L{
�B��u[��(_������h�X����ܲ��Ik����߇��B�w�&��)y���E��k�sJ��x��i���eA���Rc�1��l���qn�ߣ��q�Yno���9u���� �2�6�(L
����&r�W>~�g�F(��A!����@DUOtJ�}XO�= )�]�*%(ϰˎZ�3�`lG}�fP��L�$G�$�3�Pt
0b��O%#��ѭ�����{Oy�B��T�:ڞbd�I?<�9=��unLf��G6@�84��J��˯�UO>�x�y��Y�	U4t��vP-��Ơ5 ��颰�۞8���T�k��U�.��^B���að�����9�'Q��(�V#a���I�l�K�j����~a�m�xAST�W�%�o�5��Y?���s|D�_��J����D���)�-���R�����G_���~�2K��	��ns����y�h0+X�[������*4�B��Es� H�-�h�	�"���n����+UK�S�]��<�u������\H�����_gײ`�('����H�k�U��"',~Zy	,�zf��q妲���Ow{k)�B��L	�a��9�wp6M�(P�8�rd	��g���l}�]����, (B �[W�T�u**�[_�2�F�z�TwO�
/n�q��"��&͌�/.�.i��9{&y��C��a�ON��ѐ�0 C4�Ԉ_���2Y��9`PVE����L�P�Cu�M*`c��"�km�T�t�<��\弯�%ς�Zn��b딛�A���٨��i�Z�������}}Xh�?��͔8��2�~S1Շ�7#~A�/��H�gq��k��Â�g�O=���T�_M�ϑ\��p�ۜb I��~O8\Ȝ��!�Q��K�tg�;�{�M���~�U��ൽ6��R�|%��֡�sb�ʿeH�K�R��T�G��"	��e�s\�R��:�[?,��vu�~ub+.�E '�r��Э8�0mQQ*�@>S�_�\n(��2 -;6ߡ,��)H�Q��/���Rc{�:5�8���͑��_���`�c�f;�r\�w���˴Η2#3��c�&��H���c��˧���c$���ՃN侊\I�>�|!D8�>AYڼP�y	��ד�����0~s��cm�en!�!$�3��̎ ������sc�0:����B��T��pW@T?�����G�t�z&V�.DTv�C�y���f��f+��\�E��%OA������#g��?r2�"��h�(����>-#�қ������+�t�FI��:| U��'���J{�ϝ�>�U	bZ�&�P�j�1�%{��\@bY�G��t���+9�L"�	է�xP?���^3�\���;�|��T��fP����.�!��.kc*f#�6p�GO�~�����.�a���X4��Ն�wlq9Q8>ޢ<�3��uΎ`amm�TC+L���.Y��-�'bu���P~ �����KS�B���lfI��/�l�&��.���D��`9"0a"S{�	�Pم�B�	p�­`�4��^Bc�ʋ|H)��:����|��l|�+�����4NAԾ�/��F�@��S�C�˦ldi>�R:�k�缆~߲PV�RGZC�E�S����U�����c�6X�᜔S�'�V��ĺ���)/>�z���HaYYWA�TNe�o�=].�D�>v��O������g�1���|�ϗ���ul`p��E�q�Q�S���
'�z�@��9�/�2O3�+���vz:��@������`���Q��2e�}S-���mu�4�Κ�C<uyѪ�D!sMW���C���n��t4�
��O��3�PX
��[�	T1JPР�W���j]���'�o��*�o?�N���������Ls�����NAp��kݠ��~B�FAiI?��WX��3W��}�e= �>Of}Q�RJ�����+d��i/u1�Ki��]Q:��f04��LD2y�_` �n�1���[% Y�[~ \�bTeM�'&>�^j�h���TU�gm�p��Ş��ӝ9W}��z.B�|Ѳr5�g/��dX��p�D��#b�<T[�4-�� 7��	�m���y,�<��,�5>�c���!���1�������j��7�� F�DU��P�J^l��9�t��֨$  �2�십M~����k�лL��;Bgnf3&��DԎ1���W�\kC��j�l����?_#S���x 0��,�Z�Uk�D�`�ɩ�6� N��RM'?�K}	
���r�Y��f�n��tU���j����ا���ދ�
��zo*Y��
���b6�O��|%,��x-�����ݏ�ى0֤�!⫏�{��I��J��	����cL>( (�<��<����
U'er\���Y�V"��?��p�Q�!7�!.�#
b��Ă�7�"�H�#�D���G3��S�|�3[��On������"DՊ�k�m6�����
�����I\�U�	�v��^6��(��hF�$A��W,I�������̏	�� ����ɼ�Dw,w�y�^�Ӄ�hU�ZQ[A_���z����F}|q�����ޟ�NX���4~��ǕJOކ�8m��
g�b}�Z��M5	���I���-I�����4�]�-������l�$�9O�]�1P�#��/U���l��V&�X;��e_�+�7�Q��Y5�~C�$���7mºAF���{^DF�R/$L���LQ\�2����zl�+i�G��I�9��̟�=���TFy��v��ȱ�;����f�����'��9A�P;I����V�5o�/^�����'Q?bh�.��|V��OA����Ƣʮ�z���������s�*w��c2|�� y�;F��V��ΙZ���~d
��5�.Մ�$G��8��z�,r㸈��:��D���!%5���Ԙߐ\Ͽ�V���m�#�8��Z���/�=�u�A����e(��,:�~��a�[�G�y0�6-���_B�ש��q,�fٵ�w�֜�sѾ��O�| ��*L��F�֜�Ɋ�eIB����O�O0q�&x���5��[�au�_�
� �0ەT}y!�BYioAA�$�H	�b9n+:��[�΁h���c��B�k���g����W��~�!�*�;��qʵi�>�;.@��,�m�'�:Q�J��h!��������t�����̛}Zټ�C%+��2�����
�p��*)�E��Ԅ��*t��u�f�!��������?N��xA�$�PK, )��Q��8#5C�l@��g�G_�kK;
�4�2X�K�/���h��`<�"�b&�:����I�������g��0��	!#����ҔD��wq
�t<�Di{�(��g��f(�饟�G���X��w��;�S��P�ܳ�K$F̣�]b���y6A�U�Ƒ��������/��7ƜyUn�2�J�^}���_7Y����0��n@��Uc�����rv�	� ���%�f�̐y;KWW�`�؎&����SL�XG;��-��|↥Ǖh���X*�O
�%?%��[�*�Wo�e.e��\){gt��*V3BC ZZ�}����:N�Ӻ�!�"(�8��[��+>�|�=���|+��<,�>�O��8K�%r1i!�J�AH��MlU���n����k���J�����J?�)��
�{���f����n�9�p�)�$�F/1�	]Q�;p��5\,���k̟����!ﺥ^�C�1�����]��15[��Hr�h���&v�&i�l��,�� �+�*_4Ֆ.�����npi!��E�6ޘqL��:���������ܟ��FTCsH�\�4��@�dL$�|$b55�X�lf�=n�3&j�%���HA��g�\�L�
�2o��i�T`�\e���Ӫ�ȫ��S*��MbW�%�H ��t8ĕ+3I,��=�`�_(O.��!��s%^����J��I�L���tP����XJ��A�K۔�������X7v\ʮ���@<��#�?���xZ����~_pZ���1�<9�ɧ��9�1����q��!~�)�s&I;L�&7�ks����}�vK �*?��g�~��h�ޜ��Ė�NT�w^�' ����'�Tu�䞎��gE07Νvە�$:-��0�Q�e�����Sw��ZR�xe�S�4֊.l��B/�T�{��Y1��fǇ�*�l�6���Ҋ�#�CCv����o��a&��I_)7WD��	`�Ś�p�v���Df�����04|�r��lג�\�]~>��H�o��O8k;'�}�^�i��[�'�:A$�eh)��(�snM`[��ҙ̌�������M�f	~���U&��Gr�������H"���Thl�f�G�8G"CV�=�@ވqe0��M�5z��CՀ	��Cd/l�K�۾N+sJ�$��re�����A7�is?���O���fL1]��0�FAM�R��(=���S�"!_xh��M�}�t�yF�#��s��R����zbi���g���D��� ^�������/7K��]z(�>�Z5�_V��Z�b��3��jĝ�@X�zl�B��C���	�3B�`��*0[i�g5{�0)�zq���8�G6�N&'X>(���𫑅���[gw���b����gG��D�OVʄ\���cIq�!\�v��2 �������I}g�#�6E��m?��Y��0Z�ʬ��4��![,�Z�֨F�I���	�cm.TA�������k�iX����gN������"�);,3��Ȭ�w/_���0Zn�g2aW�c�[���2��"�d�>���g�<�w�J&��F�l,f2F��<�|�Wm˻��i^�T�h��Ͱ���^�u���:_�?�y;�����q��}-��(q.�x������z�*��ښ5�Z6�>T��Ċ��§�'��LդXe�?|���}'h�6,��;����i _O%��pv���%\ky �	�1j�3�c�j�����п�?�*�䢇0b�ҽJG�%0�S�}
��U��rᓾ47�\ɵ��9兓�j�2D���eK�ux,d34K}����?�Ս:�%}�P�t���{q�;!�%w�1����"��T��x�s^Ӊ0
���^�n}Q��:B�P�rz�ʗ�t�E���*�)聹b�ܚ�;�J~�s}���^F�ģ^�A��u�&Lk��5Y�&��!��T�Y��Y{��q����-��!D�mM�	k
�cd�'ǜP�g~��\#i�8�ǫ8�ܣUA�hJ0������E�?l��_<Jm������xx�{����}0�t}�_�4:����薂`:ǭ�&[zNmNz��c�v�"?;y��Qg�<�q7VJ�P���u��s��t-� %1 �^Z;�i1�<��- ���^c4rW��Q2i	7�ŗ�WA��E�S�\�=��i��]L�vM=)��V�M;���	��6��X=+XGHA빤�E�L��5_	�p�nX q�]��<�j��%��)���4�=s�ZўMGf�d��p\���{�c�~�����8kܖ\�L��/0�_���]�|?DZ����l���7�4|�aj���o?Hl����(�ia=����J9�O1�#t/ 4��$�!����������� j�h
}X�nO��9�DB������/���n����W��������ў��ܔ�{9�F��sٟ<V��<穢��P�T.���f!l�_2v^��eK1���P��9+6Ou��z�}���U/*�F�I�r�X�HQ��I�����RN���fU}x���w��9T\�!+�����:G�X��l|	tݝR
ѧ�W�5O�?U=�P�b4�����j�D9���X��{w��-{�����\���ɳHtXÖV�$��[y21�l��:�9[�I-m�&�)�Hf��1�	cfX�������n�E��F-r�xC�;�x �%�&���T ���ߊ��4�e�K��`�,�\g!�6��DƋ�3@<H�r�S�E���3��Vr�]������6ޡKo�7�)zm�4�Wy�|.�G��)�_J�$�u��Om��f"8����P��i�}8�@)ʑ�i�s��G�b���Z-㠒{C�3���]����5�\'8j�h���Ib�l4�1s�w����TZ����[�y��6�`��wm�I׊ӗ��Ft�"��:Ui VQ3���/�e�&ՋvC���܄��)%��vv(�>=��%�3(۶`�.�P9�L:ꋼ�)9_h����i����`��t��\k��_�%�V�a�������(���>�Z�Na�/Wgr]B2���|]�&�l��neJ�U Ph;6%�]�3�8�Z�Ҁe_[�5��i���0/-a�ļX���o�-�u�r��/)�"�M�t���R<�%�x�F�;���Y����[�����[J
�n��!%e-�+1�S�>�:ڷ��-1���Y���C9Y��Fr���;`i�H)�n1{�U���$��⒙�#ʻ�2r��O�𢶳��6���P�>�;:��)�;�]�:y��K�}}ܸXeT���{ff�RQ��f��{)�A��2h�S-�pTqM�'�-Kut+<��I��GaK���8����.���~��H �%w��h�ɮ�iפ�}9����s?^��9~0R`��5!ç���{:���T�������}Yh�'�C.�5^q���Q�x�xyO�3Mˬ.Daw����_&A쬡ʙ����LHBAq�a�W ^{�ܪi%Y��eGGAA�Jk�ˉ��I�߸ªę����FƲ����+C�vi��쯠՘���A���V��"�y(�ZD�x6H9�1��z�:���ңdO6�U���&/d����s�񈢞�e�}���ێ�������c	a,j�Q�^ϋ��ٽ���b~�}��[�%�7�-;H7����a�驃j����R�8�3���"x���ܑ�뾒p�8���n_g���TɤeP�����6�:s���9���~��[Fa�\��3^ �*��%aҝ"�S �u��P"��Tln��5��w��dw8?8b���WI���5(D�=-'� � ß�G�v���Ⱥ��-"�˶�,37��[d��'c����rA8��
L�.��=�o�sB�	��'lf�ړ׈��/q�JR��}˓A�ec���"0��1yĽ:���?a�Fw�U��)*���Ģ+H��_�#KY�=	x��r/���@Ab6�S#�"Gƨ݋�8�	�U8��a���b�:�s��Ӻ���:�������u���!?��!Q?3�I�����a�9$��F8 uF��)M�qf��g�(	LV{�se9�=�����@�=���Y|�R;	]�5)����(���m�����
���O��(�Ԍ���K[�?J�^M|*�Y�*�&fȒȳuֱ*��i���,o��i��SyɧLZ_��d-F��&91����n��DQ��ek�;&~�K�/��}����rU�c�DY�w��0N#��0��t�zo���=�y�2d���b��;�PH�2\�7�	G��Q��Y)������#�#���޲8��>ѧZ[���Ӆ�	��|�~u�o�N��`
��j�k�	6}��T�m9D�8�8�7lA0	֟���=�l"�%$Tq��J��k��&O@���
!�^��[�	>r	2c���p��k<~�Ƒ�T ��<@l*��|��i�F��ۋ1�f.��2
��%Q��r���֠c���Y%�+��r�\��"g�Gf߂�2�}�#p��Ym�P ؠ���C泺S2��vA`�	m�B���h�q���%;��uV�j�Z<����Wc��>;�}u����>@]�mgդE*l�Hj�q?	8�2w;��G��FM����c�6��U�� �1rjި��hL?�2p �Aԭ�O��!<��{�}�C�v�
�N��E��
�7�2�Jy��'Ru��t�F�}yu�m+);�s���G�-���et3m����F:��/��@lbN��t�~�I�H�<vnC�����M� ��#B�bkċ>L��<��A��"S���,�J�2x��ņ�p@]�L䩾���L�`�eztv�@�����G�Е�_D��"PH��8��h�]iL��`�A^~�d������,s(y��P�2p!z�5Տ)�,�K)��(�`�$	掶+�iJ� x�u��	נ�w^TGu�9��Z_#��\���sW�l��&<-�t��vuї��t�6��Y��b;���;�^4_�����<�p����CfF�_a��Q�o,�J�
�+I�^5������T�zO
��O-����ţB�Gѫ�TSn�iJ=���ZN�8���X�Uh���+|Ɋ�`�,��du�6
�w����6}���f��lsH���싰85*�FGdk�����O��.��u{�D��9��LJ��y/;��4����X�9�?�ԅ�+Wq���$��f���E�8�64���d�8E��J���o��Gaq�5+�E82+��"��ӧ��٠)}��ꊽEČ���] G"�Y ʋ y@d��.��N#I�ʇy��02UE����k���=�0��΢�^������c◉s<��C��K`�����~`��޺dg�
���@} N���Ҧ4��U&�d��şp[G���p����.u�=���n��T�#��~��淾	s���c��^�E�Y
2��k�W[R��0+�3�0�v�fZ���lH��K]@�b�ƥUղ��՗���͵?�?�v
�:����JC}r	P?���!ZV��Ƃ�US������.S�ّe����r�rpF�G/f�DpQ���kQZk�W���hQ������Q�/�$����b�Ԅ����o�^�h՚��DB��JU3ܫ]�i^s<vk
~H�]g>�K�ſ7�T��ś�L�k^����$%���Wt� �|� ��󩱟����:F��w��;��7�<Ga���0x��m"��#`R�����L�>Ea2�E��x���鷝{V��2�J��0戨/����|�'�� ��e��27	Θ��x�\����z�h�fF�t�FĶH�JC� �nq��]d��9���z��L$�C���z���d�5<5K�dԾ󷹏����Y�p|��7��~c���E�YPK/q��aķ��1@��&,�`l(Fi_���^uN�vg�xIJM�b�d>�*V7�����)1y��~@��M���V�e	��PF4�Ѵ�u���&t��.e�W��Do���AE��ȡ�"X�G�/vFT��0�A��9}�鏽�$�G��W/�l��;��E�q{N�4�.3�ѻK3%,h�����TPcؖ����U�*8�M	��
��L�bd�|xxS%��J��y�U��8�	9���R�������;�sm���?�9mg��Ӳg����0�Bqw�r�� !
Sj��\ ��7�'�G[?�C�����	�x`�YC��K�YM�L�1�$	CL��da��l'����·j�@+��ު����/f=��YV{�Y��r���_C쮤��(�79:-JJ��0�m\���)�RMb� c��t���1�~}J�R�����?�$s�&��S<-5,�QŚ![�\��<|�7%�#9I�'::��ݿ| [QY��*�gQ�R���k��CW(9�f�0ro�aևv8Fla"�kƴ��O�"$�vA�u؏���<k9 �.�O�iS,�Q�����	�H�*�{����k�z�y XC� /M�n����O��io���Qi^��.��"��I�:�����?���!M�?)`�|z˴��9�LD	�.S�mXH��N�`��|˾�oD�$�awY�Q����E�|�~��2��������_z���t���MW�8�e�q�u�������#m��s�
�y�}n�s9c [�^�{�AMN�����Dd?	��{��="w�פH�D.Դ�B0J�:G7b���6i���y(���;rKpw^�h��t����x����Y�s#H贄�}C�SkB���M��3^���t��	mm�'�E������=5�F���W1�/�����D����vÀ��+�'�D=z���Fsz$�](�e$�4���Ĩ{��#�&|���G/����ue5�k-T�{ٳ�u#at))H��5���p�).�w�G"�j/�-��.E�V�u�������������7��*Ȋ]aT�w^�d���+�a92>��g�Ur��6	�amq��)F1r�W���������7OU�5�w&KpjOtτ{J7:��H��HL�����G�їb��d֝s��Ք�f
�B��i@ϗŠ-{q��3�T�~�y�6���>�
�;
(�Iӱ��f�����	dP�Wi��97k��\�G�Hc�����Ŷ�hF��w��ET������~S�q@ﺙ��&UM�y�?Bh�� ����Rv7Y#Idgi;��Ob��/̃ޅ�]�޺�ʮV�1��N_������O��C.�ƻ26����j����N�Ű]}�@�Ο�,;���)����� a�!_@�/����-�6m��0ұ�����6s���8����syӘ��:���0Sl�쒃��s0�O��g�'�rw�yԠ��2�^j��w'bg��� �g�w��[d@���|�#g+�r�Q�E�����3p�a6��& 7\��էHe��]����!����̡��)m����7���.��� ��G�/�v4����0�~�F��X>&�4��0p�Y���o�ѿs�cz]��0�`�TY�K���Z]�a�� ����㞙a]�D�,��1/D|��&��O���&칍"�%E�N<V���7/F�� A�LJ�pi�i7]	�[u²(2��(��̦=�� l���я�'#��"I���x+��yu3wS������͍!���f���l��4�����u8�U��a�?:�3��d��ٔ~	G[���0k��V���ÊdXy�2Ny�W��Z���%�zp[����g�Α�:�5��Dk��q������Iv��/�!-�^i��1PK\��+x%:��sa3�L����L�Z9��qR�.�`����_q����ģd�[��Ӡ5lc�f-��Ք�7�o�VU�#�1x	C�|'�CK֟�w:`�n�I�a�k�ٔ��L�d����.�t7�� �G��LQ��j#ӽ�����}��w5z�~���Hb3o%2+ 8��ٰ��~�����gt���x�j˪�TΕ�����o��d�^��WC�o�#�7?f�x�0۱��A!�p����;�N���>�p�pV��Yj:Qs9^�?�F�x��$��"������:�/�ZX��BrM��K˻�{r��@bp�zh[4x��m���]dڝB�Za�!���P�ʆ\��0i�6?�������U�_��9��r�� #�,�K/�)g�����L���{�Dcj�K�϶R&J�	��W��M��o��+�䰪¼m5��@AF L�a��X�4.��HN�J�k� ��]��v��,�0�����c�ж���[�h�7�m2�G��,Q�x�����6�$*'��"�Z�8� Hj�iAN= �%����<^P���pU#�u� ��ϴ����h���nl�׊��dƯ�a\�ɧ	>v?k�W`k��\�J\O8,���S�dxHT>C>d���N@g���:9��%�G�1~MUy������uႇ�|3f׼�t�+@��+.��o;���j��)2��ק����(�z��%�t��/x�T��
�M{`M^5��.�ׄa1뚀M��J �;F��-��Hi��x�F(�ꞪaD�eL?$�5�p���[8�f�}U�ELX�!ѷc�(�б�'�	�2u���ϐL=覕���ҵ^�>D�Ϧ�*��!�d�%5d�$4����i�V.A�����DO
�5;��;�X�d�&9�%����)qd;��X�7�Ů[����T n(kT�����=L8;QR0{�>kjd��۹,̻Э�$�`&�����0�´�pVn=��f�rj�������dj���=�ӓl���Z����c�nM!���MJoEJZ�@?RM����;gRq�/ ]�c�/�ps�j>��oE.�~:���7����X^]���Yʬ������4���kq��d�W(��g7d!�˚?����64��{������:��B���kf ϣq�����9[�����<3!�K��@��W�Ͻ���I�t�e(�� �>�G|y�!�n�"u��*?P�
���Ku��~�S;m�\3���m�E�l����6+S0�Q5W�3��y�ǧ�����~��8����qy�C�)~��qO�|^���������*��3����EE�6_Q�kB�<�?0��7�0. J钋L�*$���kF��l҅�&��^U;l��|RҰ��6���bA�3�oZQ�-��c��N\o��^�(�oA[
Cm���8�p���ss�U5��S�':?f°H�mI���ş�*K~�u� i�"(*1x�c�����#mm�n��vf������Rl~���"_D��4����vQ����*�]���Oo�;s�����4DϋoA�5���~��PZ�c=�Q�D�`�C�o?�1������i��L4iGa���dʴ`[�;�͗  1��+-����t_�X��Fl[;-�f������P�Z �Z�aBA��/X ��]B%rKEV�۠��k���� <ln��/uZ]%rR�_��9�\53����Y�_2n�ȨM*�?dU���r�?�ş'��I�P���nև�@�a��Yu����]2�b�ؘ8p��9ܬ�ld�\�6��{7&ɎNNml�7�ş���gn��P\�C��
�v�������vr�r��V�9��C�Ox$���.)?lrW�e�D3��=5�
�[�\�l�+����l쭙Ey��!������j8��v��P�̲�L�#c7���1���9�A�(���LkTv���mC�<�ƶ2l�P���#�?w�(D@�P�����Q�`�/�a)�*�$�	" ����cI�(�2��3�T�_��A��h2�/�U���Mo��PKu�Is��6�.e�s��<��t���Tg�d�r��.�JI�ސ?a0[�S x7�*�o�V�>�AgS�<B��j��p#�^?~Ri94¡�D�3�_��Y�u<���e��	���)�������kBD�ŝ�U�Q���:��)�)�` �e��g9�*ѭ������2 �w���Z�#�7���XYn��:�Glo������6����̃���w��1��@c�L��"	�<t����ZW�b��[���h��G�X�Ҕv���ٿ����S]�r�<��D����~'< D���Z��=���8�}�@�Ќg���M{�?��*h-q&�2�G� �Ԭ��ƙ��
W�g�w˓���7ٰ�P1��H91|ӆ���omjc��[���6g@f��,L��r9�|Ӻ�D���~r���趉� �A��������������0(�$l��k*y����}����-qM�O���%J?,��<ͤ/����b����S֎�
2�k�^� y�|��˪k ��b`T=�Cr��Cp��el�<&�m�a���֣4�f�����{�rͷo��-�`U�Ak#�坩ٵp�˴"2+���d��g�j�r�B�ōW��r��/�l>�4�w� ��W��Z��<�RO�:`��٣�]Q^d˓�������R�9��$ ����� �үAcT氮<y���+[u%x���U�P�v��eu���X���3iǊ�&$�7wߊҼ�|-\8�&"�T�+�Wɨ�%��?�MT?��6��*cG�c�-�W)����I��[�JaO���<��Q���%��������l�������ʖ]��H��Jйz�8I=�,��'�߃�V�z�gdmgg�����*]$�Ы	h1�s�z��.I'�/��*d&�}y>s�k1#�����c��/	i=d�?#��=������6�%�VJ`���:��'W�X�'������!�]��#$0T���	�H��)���:E��TO��!2w����M��Z�MˎM�d�x<0�*���͹�t�7�X�#C����y���6S7?=j!��o�(J� ��aB�5�&MI�8�'��d�;�$��$�=��g,�t^m�����3ĒW`1����kN���	9�n��e�haB|s���8�a9 tB���0�'�%^[��խ����|yk!���
��eң��uZ�z��8>@(r��4f����L#i�	���W�%<�ed#���~��c��@s�SD���&����U�l_ۊ���Q����m]ZWfi�8w��*�����u9��-��:^ё����w��o��1���h8ʽ>�I2�II���;X���5���/��R�#-e+G�ǔD�#x^ o�hw�����K��� h�q�?���DI2�T�˜�I�G7��S�F�֧��J��B���H�x]������%�W�)�h���?���! � ����`( ���C���a�I��VQ�����4ZT��6=X�2$��g��b��WߎoYƗT�%jb�W�Ё�_
k�B��QqS�-S"���e��xe�^���"$�$[�i�I�u�q���R.�T��`ߕ"�X�+ˮ�wQާf}��O��
qB^�w	��RY��V�_7	ݱ����ӫR��d�,�ݡ����$�^/<D�J��)u[&����5���i��@D�!Ƶ!F9�D1v�o5pJ,:P`�����B�Y�Ca�P�>"�G��<G����?��X����T�y�m��ȱ2_4�n����V_�Ծ#[0�N��~ E��[�U�˅� ר[=���S0R7���C}x��!#� �������?�Q�[]9� �N�4�;�TWƎd�4,�`C�O���,� <�[Ҧ���N�Ɨ�t���.�������.b>ǌV���`�N�F&�rX�a+�>�c��{�_��p .�˝��ŋ�6:��F.��]���Iu�Jg>W� 3Fbx���@Z��P�f�S��x�������[�����cs���b�d�$��T/1����oD�����9F�W�W�u�/ҫ�ۥ|g���I7�>�Y�e{�4�[/���a��b��5� ݱδ��,ٗ��䣒��S�M+���Ť��ɦ�(r��S����A!��2�;��?UΑ�HEB��游7�gX3ܟA�tȠ8��#y���N�,�5PrA��W � �۝P��/eqg�q��a[��iuH'M/�8%�HD;u�K�`c&�0wg�HEW��_Ľi�+����y���[!�9�&6���<���]P�U��@�lT�ƪ�W5Q>�Y��)t`�7�mdT9FWH��*�Ͻ��9����b�۷͵�z��+���X`��� ���>HK�P�%P�s��%�U�t�'	���l����-jA8_9B-c�Vv�Pd42���[�c����C��e3��q::�h/(V����R�e-'���C�g(Ҿo�9�b�?��f�Or:�c|0��rak�#�0��#�c����e����]G�����ʗr����99������[N�M^۝�SAhE��a�{�Dw5"�(��e��\�+ѽiQN���DJ�� �P�<�����V<��,d]K�y����匶��>H��>�?(�0wi��S������.а[Xy�WX��5{LrL"oZ_�X�!K`�Į��4����;�?���c�k@ )���Kl��d���J�d��$P���6����Ϩ w��
�xPe2�J��F l�;+ÁMf\zڟ�V-��Z�t�r��/h5�E@ A�+8H��:~�v�%̃ E���2]���Y�u��N��?aظO��Q���&�� \w�����=��#uW��HlܑO�	S�W�>2�Z '-�pg w{� ��EqZ��w��K@�� ��Mo��Q�Iǽ�¤>,n��/6�pRD��[�O<��[a�ѩ���k^���i����ʾ����ےz�"[��V� /�X=U�K�KY�/bR:R�ӍV��eA�ܟ�ȱ�,�{���������S��\e�:J
�Ux�p#]����G�6p�7{]�n����(;�m~,@�17s�t�o.k���?M���3�k��.ct(�4�5����eh���l�*�M1�;���}Ʃ�	b�Z1�fF�w��^�����F1$�ا��8��yjW��DU-5BK�c����k�w��{K�w�FG�;��c�fG�֛ס��#+9P�$i�Y*@����k�O��M
.�yqW���~6@���0[�*����B[Ȳ�v����6�%ͻ���lo֚���T])�.���Yۖ��fi�|�̉�z%���iS�4�����;����v�� %���ۣ13f
]�!!/�q/E�w|7���K7�Yu�H	ʃPlnS�ϝ��&��V2�Ӌ;��eJ�0:!Q�4&�B��<Y�l��ݯ�v����x&�m<���q��I���P�Z	̬x	+y�O�>��	(Y�{��y0���7�ae�����A�t8(���ͳJ�/`�R=��10��"%ew��S�K*ߨ���]��v�G�dAB���=Z'�������(YV�$p6�n.3ϣh<daZLc/~
OUK�0��Tl"�ʏ����#�6�p�����#��YȜ�m��Ph>1z(�a���'!0�nd��D�-_!f��Q�n�C��ޝ�Vً&RT~�t�35	�'D���Y�[n��.��d�.��(=�ҋ~��S�6��x4���U~�N�[��<��n���b��P��������Y�뿷F1����Y ��d �$����&g	68l�Y�J��*����yDε(`���o�=�f0�������nm�E�����1�pj�+�}2[Y"bhdr�8b�5oO-c;���D��/C��S$8�JV��q�Oz����d��F��&U��f���h62t�r��ǤG��W�̐��C��srE�P6�|�4�h�R�Jr�O �r&?9�%�a�*��ڒ�ꭔ�O�-�ɚ�[L%�i���Vf		A���>Ʊ�y�<��02�$��y�)E�#	���	��s��;k�����%%��u���[�HHH���w�6Z����˵H�6��"y�Z}������
�BLL����zWEK�ji�#T�P�2�{Q��˄��=��.��a�������8K�C�hP_	��ň��Y4ÆB�L�e�l����e��q�@/����-C�4P�7i��I�GjI���N��_@�r~	�2�=.�(x�XG�t��� ��=����i�C��� �D�2�ʓ/\�cI���rƮ �?7��׭z�[�����ZijL�8'm�����I{�,̷���(˚� ���d5D]��ێD5��}u���c!N=��ß8ְtTp���@�s�uL�^{=�����}	?����I bG=N�u��DI�Su2��� +Y@��}��U�����Cc��`I���Wܭ���=>�-$INF.Λ�WR'����gcF�:�m��L�B�=\nm�žK�S,�;��K������+���3�@P1o��z)�(Y���3P��.�+į�bX�SZ/4�8�F�~�"׆)�I&���f�l��$��!:��C�/2��y���!����.�����$�l�-���M�쁑P1WrM�����h��	H�
��R���$H��)��{$/Ά��;y�{�p�=8'0�xY¬�oU��F��W2^���B?{2eh�#�p�rS4k.Z�X� ~�х`���v���g�:��#����d�.:����tI�.	ZeA�3j%��L�(��z�N�@D��b@����&��	P�Jzw��!qQ�����.S��%EG �!}M��C�6U�;1������r-�N�^�����R�g���O�e��q�T��s���Z��k�v��4's)@-�#��K��g)�q�?�����$}�4u�JB<�<��c�C�P� �4$�����(�;`��>~�w�x�m*����x�n#�t/ 8���3�
�
���ޕ�ޛ�CHk�wa(�c��\�y������L��ePF���wq����f�����ݱ��I���_�����������Iܛ#�{E��_���c��J��=���`a=��W���������`�<�rМf����,�4��j��6�Ȥ��C��7y�z��vʂ�"���c�nS��El�-�Q��t�5�F�)Wk��W/�Qj:.f�CS=�Ŀ �����d?�:F�̆��>�8Э]�$����+������WL�-D��=u=#y�ٶ��j���/t��.�1�?U'�Z�����-Ռ�7}_���xN�\b��d�4R��f0Ww G� 4�{ 3{
�F> X�ѯ�ny��?�^�Y�V)�Q=`
pͫ�D��t4���mY���I��O��ש�b�y�ک~�����i���N��-Ln���!���K|P����}N&
��in�@f����!����p�Cvpjiv��������˯3P�;� �)�E�}�̄"q�>o�ۉ �`%<�ϧS���#�٥F`��C�u^�D�G�æߓ/�\�W8��;�/~Axۉ����M�k�f�֜��ZTF������v��_�r�'�����G`�k�7��T%b�^kH������"�\'#^(сϜH��g��Z��r�1(j�ە�ٴ�8��7��.ʐ&�7Z(�5]+�2*=�a9�>�͌:��~X��#H\4��Ԁ����om;����9l���mp#3XX�WI�Cny��
��j�[���e����_�*��pV�e��""��=/vC'ZP��t�\�q'��g���C�F}jb�죹^�kK+�T|��W�'�o� �\� E(���|"1�����(*?�=NN,�Tĵ(�8�aб�]?L~e�O�b�ŀ���p�SiY��
����|ʲ;4��`��9~�nq�O=��F.��$=�B�Y�9(�>릙{�eUL$�3�<�S~�V�%
9Aኮ$� � y���^��<☔����5jJO�J.L����
�NS�Q{mܧL����\!�<�Y�'	�u�Q!7��Y�Zori��4�Q�*&���Ɓ���H�^,�꾕Z�	L,�2#Z��bC�i�(y�)�ڿ�?	J�%�(����K����3����9�t�I���9jE6�E�� �igw{��?�`C��v�OD5;�r�G���j>bl3C�oa���d<���_5�r�4��|�DRYS�*���5�|�SB�^�����w��#?L�T���*v��t����ˁ�־똄��I�ag/���E��ٿ�g P��#��؆5}EX�s,�(�C!���F�@�J����_/��Nר
�A�d��(%0~�R�L�Es�����Æ��@Jz�����4r�tu"�Z�u��3����}l���\��!a�N6�ͅ�" ��5��!����SW���lsU����?P}���)]v���aE�q����0&�
�Ú[u8Ш���!A���]�0��;������J%W��1	<�,)ö@1�H�`�XK�� ��0����3���hH���*��4�Dç���t�掠�e�G�D��h���r���U�XJ�_��d��s�����ʠ�~�'���P��УΓ���r����0h�����\��A4�:a�US�R(���vPF0:�q|�9'�4��Z
]|�K�Χ��6�Z$��4�Kn�J�l���iv1���^��w�g��O�(�p3��� �s�����נ�}q��d���i�k�9+>����׳�MҎ?k�?�҉��:5/�T��K�oKd�@����C��/pp2AO��4���/���ё����t�~ۛ�{N��᰽��-s���3;�����������EO}Sf��/��Q�:���`
|��n
_�n��ȩ�4��;�ȧc&�;aT��&n����	_�F���4�<@�O��lGJ�KWG5��5iA�&u�
r���`���ׄ_}�qd�J�~�˭����8n�|oA^$r�<y�Y 7\��`����XQ����Y�G�%��o�<�����L�����|��%�^����������� )�?۶a���6���^�\x�"s=��(�a�0Q� 0x{j�w���~W݋����Cf�4����P�[&�$�a`�}B"�D�q����v�1W��<�J5����/�����-	��b�-Ĥ���$�
s�USߑ<H}y�ҟ:�-�O��!u��.vC�Ʒ�T��i�XƱQؙ��So��dx}�JtIF��z�4{1���F鄪�g2bzBV4��3��з �Ń�~�lΓ���"�/�pH[�Y�2�{��&�lp|�zK�H�ߜ��I �$��c�*��-�r��c��/(n��ֻn����T�)�E�e���8���;���)@Lm���GM�� ��5d��q���q��s�ߥ%,l�}@�aF3�Po�1s�<I��F�c5��↢������k�c,�Z巄�e٫.�W��`C0��i9
W�6�{W_~�e{�/Ld�
*^�:�����/�]��0Q�yB�����^)/��R�f3��+t�i��#'�!]���yr��-_z���8�zbCYA��N�0��x���z��񨲚8���#�������ި>`J�z����H��o;��3��{XOK6= H��]�D.������4\
�)N� bؼ*ĎN+�>�7� �J�J�갔����y�#�M��8��z؏γ��bMZ5p�|G�k\�o��O`,7#^&��v��	�p2��b6�&�Q:�N�U7�ů1�Z�4b"J_7����b�F����>��'�~��<�0�<�a�ړ�`�߯�#�o��f^�b'�Ir|��'3?��F�Z�|��F�g�V�/Ω!�@��rp?f"B����+��5�@+:�^A���Ḇ�@Lo�d"��L����7@<��y.^��-�7��hLN@ah�Y�"m�y�y�UC����(�-1� M��CV��HS��kBm�6��p�^�������6k����'�H'��5��L����|Ӊ	ҹ\^˗'������@w]���d��!����#yq��?��xF&�&ᤇ�WQ�A_�Ѽ��(��j���r	�?��V��O�{�9��a�H�ך/�@|�N�5@PWI��r\K.M��;�>#��?���4դΘ����ɂk8�
��.��������eC�U <3Df$�eZ����@��T����6IP?kn�	Ǚ���ʴ�F�,n��ǥ������}TzɊ�yGĨ���t�o��g�*�$ݶ���q���������k�(�
�ȧ���ɬP��rkn��آ��Y�
P|	h��v��E��ϗL��K�l��#�h��Дҕ���`l{6��g5���)������š,]��I�p�#�ӄ4�oaz�m#%G������,*���?�I��jQ��,�"��8����
P��M�>����-�ԕ�T�u����tJi��To��ގ�(�\�"�##�!��J{o��m�Y�G�g?�f&W�4��LH�K����2�G�m�|��9p��f����_ 0P9_Pl�Ƹg���`���<���kH�獔�5�YHʟ�$�C6ʠL6�0V�`�0%��hôJ-;"�=�������D�r$����]-7+6����S���5��O�sI���*p�b�U���q�;�9�n�c�SD�RDi�']���g�8�n�G|�|��eay�sIԬ
:h�&%����y��_��=\8�.���/8g�o�ٕ8���H�=�,�Ux.��Q�%ߝ!��x)=E�v���}�ק��N�9�0���oȀ�B����;0(����V�X�	�7ۃ�H���\��@��L$�۩��ƟO�����6`DT�Tef�H.��1�r�Z;�� V��i�[����V$��B��݁+�E�G"�Imn5�[(o��Ym��k���-,$�N��O��Q���fv���oJ���C�}��d��k���5WS����8ծ��䵅�g;�#⛡����~ɥQ�
���%č T}���t� y��E�>�e�[�>X�7Ey%����]�e>
^臾�o%A~o\<Y6���g�� ��.N��D����J�8q�6���_c�Zj�j�O�G8�dC�㯤�<(UC�#�;/������S��CF�WI�j���_A"ygw��HwY�&�s+t���P�^�p�Ҡ��E/�ˢ���t=���5���3Q��j�+��o͔"��z�u�B�yB%���BN����e�e�k��H3��w(<\���ӽ,i�}�d�~(��U�E���Iq}�@HK;�Ֆ?/ѐ�1T����;���I�Q�ƀ!����O�6e�!�%�B��ƝZ5:�v�G��p�Ee����P6�$�f�j�"�T$���}�@[���J�:�T�̆���Wv���ɡu%�R�
=��;�\`|�SRO�'l�`>����U��"{b=�L��l �c� ��SDP~|~n�R�
|"|���dz)b�v�C�&���Z�;|7= �vΜ6�\��-݂QI"�I�b|�"Y(��II�%L��C���J�ź�9��S������*QLǉ���iS?B��#V`�����|Z�^�-Y��6�e�p����<	U��5���R�m�_�̯�7}��4�c5AJ�t�d���0��u�A}B��R�҂/���E���S��ci6U�R�zU��Е��W�'C���GfN�4
���ϸ�����@qY2�VGN˧�H�X�Q��N��wg&h��Gcȃa�i㵷�Yn��[d�S+�OlN�y�DI��ۢ{#�����6T�}�E�ǉ0v@Y�F��@{j�a[?Y�|�E�XOl�9�y�E	:6�*�A'���������9��^/���ћM8�Y|�f��<ll��7�)�{>��)�	J�<�w9�Y	h�E֕oL��p�����8_
p���T�o����ʕ�����<NVĠ0<�ţ��w����6>I�31ӯ�G'X&Fg�(���������z
sd�5�h��ܦ�	M�ĀR(e?Pb	�������7Pt&��b��L���Lzh���
l���aVSZ��\1_*<�ָ�z_>�V`�eD�g��>-�=#��dO����)&Cї#<�Y����4�|@�L�T�L޲�L�,�mjwd9W���bJ���JY|=c��/Bx{�
�a��w����R��qS-MX�)�٭ӼE����=�����Ջ=�H�f��Ŗ�p�u"����j��f既���]��G�iB%���WXH]�49�pU��6��v��}��C��Z]�� ƍAm���$�+Ԕ�\�\f(�L.m�ޒ+(��Ԛ�%�^8�L�i�#��ʗ	}<r�p�Q%˭3�ѡS�:�����p��h�ĿBL1l���U'|cUqQ`GF�F��UJ�;�H}�YA$!W�ʓ�<7�Y�S~���u
��j�p�>s�w���M�6�������ԗ��b�V`�e;G��CL��[ǔ9?����g�h;"�a��dG^�t+�"P���*����b���#	/DKw��o�Ob�[��Lm+X�SN#�|��<��.s��Y(&cG��H�3�	L��x�+dy���M聶w�A�����uR}r�c����1�[��k�-��J�;U�[M� s���zp�!@<s�,�����~��97��K%��U�,��x��B�WL�P�J�6��;{nC��7j{�<�( �'�w�Y���-j
o�*�D�ٞ#.+C͡����/��n�G+׶A��k�Oj�VM��d��Hj���b����١2t)���y���%��fƑ���@��K����lg%�,Aep�P;1=E�?GY�XCͩ���ϕ=�;S�)T�-҃�&�m�#?�u��G�%�$6q#�r��G�[f'Љ�?K�FsuN l�d�!Oz/>�p�M`a����b�yM)Sj6� 5�`<6�P"�M���%9��RmT#������2ӗ6ruS�4[;���^��k�Jh�$]JëK�nbt�����B�G���O(bb��S�R(�:獎��d�ڹ�
jh(��g��}Y+͸]N��eѲ1�ݦ��
���,���R�#�=V����;��o�1a6c���x%��qa��/y���R�5EXB�Rʻe��j�m���X��+���&q+��y��:�OL?��XM�Ю��KP�S���Ϫ-OK/�OaA,9��6>�3׷��U�n��˨���`NK��a^����d ��o�_���Z]�'����yh�|�h2`Ƀ����z�<��� ���Qi��fyL"�fUOG���]�Q�;����㮤�:��#!j��yH�˥�{#�#9�蓮p7�h��@K����!���$���j~8�1y�'��S�v��p������sN�?�8�92r��� %����J�x�s8�s�T�z����ޗ] (�Z8%	�*(\3�>	0��>����n<���\����ݖ��т��`�X����D�j��"[�׏�Z��v����J���)m�`�;����̜v?����J�]���K��GX��<��%K5?E�F�t ��%��<%읆�Ʈ�!$=��8�nF�?{���Kd�"P�@��_-iC��+*���]�O�I|_3�p���H�o�(J���w�f�6���۱�o�ȶ�8�g��g'�^� l~�A$��{^kTen�1�u���A�_2T��dQV::��X]A�����0*���b@�6p-�M��<�?��
ْ�Xݐ�S��)�8>d�4�g�LK:{B��#�N`lW�ѫ�@�i2�_�m]^# �Kr�
P�cmlX���1�d*���"qM,����X/�=�*ƭ�`�	Ml�@,���`�a`k
��מ+|D2[^�x�(e�9�3
�&v+ڷ��Ϧמ���r���[y���k}�%}�C����6e2u)L��P<?K�>�(���X����;t7s�Q�i@��VI�6N����D��G"p��)�00ޢ�B��f5u��r0�X��7��*��c?�/x��]J��uKMP.b�4��ˈ&ZUk��\s RqbB�s]�;�I����aF�4��Դ,�B��a	 �����u���I�����'@Պ���m��R4Y�ua�A\g`�=����X�0X޸C�*n1�M �����:9צ���P�]g�BD]��=� ����A|��w>���a_7��t�Q[a[0�mB�!ʤ��ѓ�/M����my]���i�z5|��}L�Sΐ;-��+��_� 1��hlj����v��í�`cC�#r�lʡ!_�K�ck��%����G�7�
Lc1̰����v�L:]�U�Ԧs��G�4�1kC<���yE|S`���2f%ʃ@�����f��d�����煓 <G�c3����"��]
֩ر)�k�1V��2Q5�D��k#��2/���t�����{��^0�)��;�;Q�E\r����ڜ`��Ͱ�}��yu�hA�c�ʣ+dcE������{n��Su�cM���v�l���Dо�.�A��k	��q��X���v�TF89�P���0�u��҉j�Bc_��br֣~��x��Ѫ�[�V�gagt�	���n�v8ĥ���w/x�b�qN���[Jl��3����?-���c�TEJy`�R�M��̳X��#d��˺:���tN��J��vL
�鏢=쭌BKe��v��r�U� �M�򻵈����;t�&��'��@��U/e�~�ݚG؞E���C��S�5�6�,�}��o	N�p����ͦ+@�y�}��;	���gwP��y��e����"��;e|���!�MxP�ټi�S�J��4�;"U?��@|��'6�c%�n�k��Ɔ
���h�Lt��jFP���n�����XJ���v�k)�(qID���*��cm2hV\�H�˷���ic MA7V��'��PZ�~O�?�e�8��&�^G��'�����/<�P<)���RkY�i�2�n{B4wG�K4�σ�x3 <m�3%���*��C�l N�<v`�^�d������_����Gu�掴d�7���fS����L,���:��Z��~x%ES�Ƴw�q�����(�z�,�:���bP�d���j�3�p�h+��
{���#�l�9�W%���~�:����Xm��p�!�Y�Ǎ�7��;���N������z���H���k�_�˰�"�n���=�񀬐�|ݵ#ɩͭӚ�|��8������)4ެ7PF.l;4��	M�����oB�KY�ٌZ�A��.c=u<;�A�*���D�e�C����eH:���0}YV
|�)�����:X��{P�����~38At]�\��������4b�7C��X�N)����� nW�jyf�}'��ָ`��	A^G��3��C����f~�iO�����@G�i��P�֯�#�0
m��#I1�����~��������`��.�Q/���_ �s+�.��{#�%��C��*�3ǷB�T|1T�p���v��8�ݚA��;]�tjx���Bt�����-s��$��y�8o�3�_�%97�#=��0f�Y%4�A*�v�;�=ÿ���Wt��X"�5]핬�導]", ^$!�$��T�ф����y%��K�֊8�d�Ժ����j
$u)�+�#5n�lY�*�~��`�cK�	�T7�Vꐠ��_�����v��L�#�/�^�v#�<�/�6]7n3��-pt䇟�%�k��Y��F���@ٗ���
�d$��+R����%��6�wq{Ә��V{��j��g��x���@djtD�IZ+d��S(�A���a{������D+��|'Y1�8)���3�;�b���L���~Z,�hd	/���u3�yY�|*�Ō��yyN�}��C������S߱~���o�ad� b{�1�
�C��ym;^�ߐ\�4�{Sɢy��_�����[��l�E>��A;5u>�ߺ���-@;3[�k����?�#��J�جX�`UWŞaQ��0���gb�k������nxI�<6��j�.�	����u�ӯ1�"Tx�O���XGH:|�O��G+(�9sK��(¯j�D�>WS���wN�/d���tk�b\���m�畣���D�k`���A�>�(h<O�Uc��oP��&�PCg��C{�d6�Пt�ְ9Ѐ�Wx���G8�N��A��P�yY��iϻ��q��,�9����s�dv+�����ss��u�7��;��}#��򭣳W����xW���d��/m!o~X���9i�\N�@��X�ϟ1��ء�O�Aƈ��*P=��y(��UHG�ʽ�Zl�䂞�4�$▙�c���r߮eWe����C���9������vF;j�v\e�;U�Zu�j�)�{�GS�R&Ƅ��.�`�'�u�\sha��P�j������o�
��s��v��*�OZzn*Z�( r�_�Ц5�7�&a7�K(� ��~�OvֿI�C! �R�]��>4{���f��Xzܜ6)��Ғɲ�>��9�����O]���}R�� �lr�6<��<|�<uq��v�w�SD)���x%�Ǹ�ħ^�8Y��i\`��3'�0�L���Q$Z+��:|'�U
��L����/�y��AjH.�UշGn&�r��+���v�B�_���CaY ��0=~�JD���V]
3&�Uӫ��5?<	��n
��	�y]|wt�9��pv��6h���ݞ�$����|�0��C@1�1#�"E�P�WS��.b�X2ap�.U05���=�2}`]����E��")�5�^g@+�25�4.RR{>/�E#�WR}_כQT���ߏI�䠖H�\T�R
ߕ/�{��a�Z��)#��!��%�H�wGN��Qi��K�d3��0&2���Z��E��*X��H�������N����&�h:DV�|��i�Uh�Pu6�gE�JgU)Ԡ��nbš��l1�
�s-��f�=. N���[=�����<@�����R>�ږ�}���ٓS')G(���q��Qh�XT��
��\�5⧉a�\O?VUjb����mה��{�0XJQ)"���d�;RG�6�,�h�����:� �>O�0�Q�V�Y�@ac��!�V���"�_jK/�J�TY`j��!�s���ʈg�e�?�����9\�+����0�:#W����ʵ���#�͇��m��M��@� j���_2��N�,+�*p��� �D8z��!ځ�w���bm�u�X�Z{�_I�i!_ט���;\�t�ꁪP_�9�8������~�0n
>O�1Bm�����	_
j�k ר�C����'��'H?"n��]c�z���:vݨhХ�̭��)pG�+M��`�b�ƌ}ᵘ����
f� τc6�;q���}piG�΋
�.3��Ӎ,�w�����_���>�9>։�����1��]���*�[Q��7e��ec�sJ���t�|��Rv�@���t�q]�&��9��my���n��VR���C��:kn�&���ۻ��ߡ�M
lq�[�}d�f��.��ri��L:l!�Zrջ�Hۤ���*�;n]'x�j�����Y�����1R�;(L;P"'�ۺ_+��&�Y����7g�gJE{I��ɝ�m̜�)���.�����F�������NJ��|�j�|n�f�����ת@�N���j0�Mq��FO@��(��N�]�d&�*λ�PV�LZ�~���A^��G@p�nΕ��^�8g$L'�Ȱ��/﫹�1l�f����p���܏
I�oJq��%z2[�.-�]�H�t6	%k�K�v|_��BIiB����p��ژ��i��,�7[vE���H�"�P:k� l�D��-oT�.��΃<���>*6�X���AOF�9z�ێ��X�f�˅�ٮܑ_X�x`	�'��� ,vi� Å�[�肷arQ5����t3�E�(��vML��([1,j�t;T�$=Y�A��ֺ}&%��vܓ�`�����5,qi�z���#A��%��1�aQA;��dk�g�a�,����� �S�uɳ�fy��/.��5䌱�6!�z|\v�~`�H���0,l�6~!Br�z��.�}^x�g���g�\r��v(^��[���Ҝ�;�Yw%9O���7>a�`���#��_�y�ϻ�3K[;��Q�V��u;:YE��̶�霄��K�%�o��ɻq7�&�5	�JʸӤ�Q����D|��/���j�"�S�����P���ס���J�N�@�\�H��oL�L�nsL���$�YK*v��0ts��NQ )(�����s�}uB:;�	]q�
�=)�a���/p��p$��g�-��s�q�`><x�Z�@���>H�U�\��K�k�Y}^��Z|��$pz��g=G���l���/���X"r'��q�j_&�y��h!�bՐ(���]`L�yA��S��Q0���*cv:�A&���ч��q�/�9����
��ANTՇav���F��G�$�G@�0���颳q!�ѹ�V�>��8��~���p�MbJ�A~�mt�C�����a�%�0��Yy]��s��Բ%<�>�����8�VIi9G7o	��B���H���!�r������6������.�2�b���U����ǧ�k�(P}��&�c�çYB"��I��V�,F��,���I�pj�߂�Ǝ�Ӫ��6�umd�#|�C��!dF
��.&�"���!m:� {��kpǎ�6�)�EE�\��� �']4p��ȩ��cy�5b-M��:
g�K�Rc����j�����-!)�3���(����s���-�δBfq=��!��ة��``�Q$d�kX����x�xר�����yy%�l.Q��LM@ˋ�erX{�bn���d���h�+��\���D*����{�L�w���]�n�%>e}��Ky�fuQ:��!��t)\N 8.��	]��મs�pr\����O��UdC~�^����1�Z�r�2Ζ.3���Q�#hF���4Lw�z�|������ܳ��C-Η�c��zc���a���1Y�5P�+�Sz������|�����j��༻�O�=B?1؜Y
�{������'u�u�*u|U��R���2M����2aD~g���ء��"�����`�C�R�QI$��O���ݭ������Z�T����;��U��m}�:tB!�c����f�&%�Bit� �lQ_�mvv�1N�;�8��g27����/S�ٻS�W���1)�g	{#s�#�A1��r��Q�ҋ��$^u���B -7�gǝ:CI;���2��E--kDvR�h�=J�(�(=��.]��2�n�(L!���[��濐E^���֬�*��)��;��&7��h1V�*�B�w�5XI�n[Q9Ƈ񟄋k�����v�V�0\f���:d��*���w�3�����:�"[���[���;��Z�;�"duX��ۚ����B�#���g�V~���<M���*Q{�<�8��3��Gs�|��,������~��iȹ?�r�cq�S�=Y��}V���]P@�(tIɄ��L�q
h���P��˖����g��R�3���'�,�TƟ��:�8��snơ�4_�k�H �`t�?ʼ֢Eo;�kWdU�@'��r��.��1��|J/L�+qkJ&��H�;�_ֺ��1��������,�q 	�^q)�W�Oz�z��C�%��PX�fh��_���hF�lKrp�����O*�ZG4�0G/��P��l/�d��,>���U0Ӭk�Տ��w�i�WQ�y�q?��h��b�1�%��`ܰ"�I���c0Gs��8ΰM
"���s�9*�[�!H@��8��ʋ��r�/,OD�[�!#F�+����h�La8�E)�͔��(���@����@�Y��y�i&h�`Mb�]i��� ie���G�$��HR�S_�De6ڳRcaF�l�	�5����-���C-���YO�������fõ�`Pz��A���,�Zh��i2j�ym�[����]����
/���E����.���d�{"��B �����gBb@ߔ��r�K�$�G٩� !��iV��L�������Re����w3yK1�br?g;��ml$�5�Y��h�9="/{���W���rc���uJ��k���:�s\�լ^^�Igh�+#E���ŀ�5�~��^����c�2%��^�C:td$��=5����N&P5�D��8�L� ����g�LY�M=����HU'�̺�i��b�[p������+����	{�!�&9�}����^�Q�M�Paj����63MtrL�6+i$�/OO�mgR1��S�ŵ�tBz��h�P�\�����lт��}����� ���6O�(¹�蕼���}�0>d�����N�`���N���m��@t�LrWV�ޒ�r�7��p{�Ѿq���r�����9]�lJ�";�
�м���"�mq�Nt֖'��(Y���S��r��v�קZ�SϢ �1��$�pu}��S���ڻ�*�
�ut��L���m79)s���X�Y(���^f�EJ�ߍ�'�z���������=|�a��h�p���Z����{��d ��W7ɮD���i+"������x�o�QU�5�v�գ�Cn�X�΁�Z�2���޽P�d5�+@�\�@gb� ��>m���9v�z��.Cl�A�����<��l2_��������H:)Ub���&oP��(�P�(S��Q��21j�a�U���������
zp��!��L��tu��+��9,Iy�s`7�lb
g��D�v�m���t�����)�`]�F�χ�<3l㝍������J�Z��o�#~D�x�m�7Y��x��K��ۃ�G�1��60�ey��WiV�ļE��c�`���~s���A}ZM���l���2S�К�<ڗ�0[Tq��`,��\1��KN@����ji�S]��|��u��7�i���/38snY��^h�GP-;��B��^��x�$D7��v��_h��+I��ؽ}�K�}v�V&��Y1/�5���^Q�Dr�Z,��C����i'����x%݅0�5MiP1�g�U�o�� ���Z�m�z�������%"H*�h���W+ŁJ��.��O�<�_���<��YQ��ǐ ���SrE����B�F�D�b8<�@QHm��r��>VVF�C����<�g������Ԝ��sLT��>��0�X� K3�h*�0��y��Մ�h]��D��kD)���H�L��>����@U��m{%�%��T���b���Wŵ���g��Gٛ�Ċtz9�I����_n��^����GX�D�_}ļ]�k˹+ӭ"ǪȦ���o�P�Y8鿀5bI04%�Δsg:5��2یS&F3�.1q���y����߮)h���Л�j)꺔��$�]�Nʗn4X��X��|�����إ��I%�c����)��gy�6⯀ٞJ���6aO��C�4��%؏P�~���}B�'�������o�iJ�8�cb�ګO�4��! �(�]A"[c,�K�5�=�	�q�TrB�gMyR
E �R9���:}��p܂��g�2���w���$ l�)��鈅�<�d
��74�>e�*=j�aP@���6D���_ >�N��+"�A���QA.����e�q�N�j�}ٷD�J�M�Ub�#DC���i�:i�k9KW���D+�3g��.�[Y>*�/�M�/=�/� ���4QP����fN|���%�C�	e�-D������oxg�~Y�&|N�X���L�`���*$&-�'�\��	��7(�A}��/��
t�櫀���e�<�d�}%Vwy}o"������Ēշ�U�%*������ִ�M�*���>JJ,�3+Jt��V�D[�)�&|�L��Y�Q�b��[�>�@�#m��,��S5܆3W�5cs�t�;0�h�}�x��Z{�-�s�et
��L_�X���4K{+-����}����/�>�`H2�K��Ȕf�8�.��9��xDMB�Z���5���M��p�{	P=��C�(n�r��)oJ��?�Ɋo�����v*lsɂ�MS��+���Q	,�N�I�%����SZ����4f,k��ۀ�0�Dֽm	��8ݝ"�1ڡ�/��_�"O���89;Ҩ���vןǢz�����
A�k`�Æ���θ��#��zk���Փ?�/e
`��'���2mk#��r�q�z�9���^7��E�U�V�(S�_K ��H�`${��:��QY����rfFWt��'�$�����8�+��$%�HM<�o�5�Ԏ{�#a�(T��d���Q�e�قʤp�� ~�1s8I#s��������i��5l��.��-�f�c���L'�ǲ裌ʱ#��\]"����7��E�]����^Ñ,��4{C���^�b?��o��I;�9��v�y�Cd�O���ه�������/G�/yv?R�MvN�}��6�� �:}䟆��q���]��KBs�_O%�|p�j٧���%��8���B�O	#��h^�B�n�m�#9�x��P�+PU)$A��M+=w�G��S��u
_��I�������_sZG0�P�5�� JsIef��Av��G���} �u��d��T�+7'��8y��d6p��9��}���9����}t����HZd�={w8%S!�����ȑ�����.ME���z�3�Ih�z��7{΄�c�Y��������Z$]����&S�4V/�ot鯢���R�q���n�A\��s_��$�����3#�)��em�)U�k�t�Z��,�{�eZz��H~	�Q�p�?F�[��aܡ��y��o��r@b<;.I��A���GX�0�u"��/�.��Bf�b	"ߕ�sx�"j���G?�"A���l�n�N�,E���ϓiI)d�ʀL�<��<ŉ���:F�<:Z%h�
�mb���4\T��Þ���B�7y�3E�����꾡!Ӆ�Mt�pɻ����3E�	Yy18?����iDq���	�N��ݞ��"E�5lw��s3�c�7x������(o�>�8Py(��a	��J��2����#�܍J��m��D}v�Z�)t��n�q#��~�b{\�"H�Q��#u^Xo1�vf�x��A�_������n���̐
c�'wY06%m-O��1��@{ӇD����X��7<&}HK�&-�1pa��W��W�骖����4�6]��a��y���`��*���bS� Q�F���Ƣ�	y�E��w ���_z��G��5B�]�c�D�!n�p���]s)�۟����lxK%OXP�`hVT�f��h��{N��D��绉���b]E삄9ձA�����_:��q�����S~�H<)&OӦ���Xݮ��5	����g�Y�6�67nF�D��� �c�&��� �F�	�0�C���u{}�Q~Iujz�ň��m����\���&;ilS�h�_���U�y�8v�W�;g�+��ڵ-b�dx��iBR�@��H&�'�۬����M��p3�L�P�0u�C���5B�۞:��.�2u3�9ų�M닭�*����V>vy}��v��_t���c�E��&W��Y�"�(�p��D�%�!5=g��'m���
N���ʪ�Q�Ɠ��ԍ�{���ʄ5�_�S@��'4��N�F>hu���Y:�Zs"������m��#�:-~�ϣi+�a\/nO87�a��ɜŽ�ů)( �?�l�[���ѧx�&�����	[PI�E�&W�����k9A���6�2�+�ޒ�w`�T��^p�S�q�>��{�qU�����������e�ej���~H�<4s����z�Xdӹ'�^�����'E��I�SL������Ѻj9%�����\#$�A��\T.�ե#q�U�^����R�<R(ֳh���r�9�͑ E����`U�\T�d�)�A�o�w��Ls���Rc�<�ca�
ɳ�#���n�	^���ö���W�IrDv�=��\�H�Ƭ�NN� !� ��@�JTZIm��0ц#��,��j�~N�(�k��&�E��=W��F��ף��z4*�Q8�^�"��Xj��K��K��x��e�~��^
��%z��]G��n}`�T1A�l��yw�.��\�W\8#*��
��:���"�#�nI�_~Q�5�K�v�6�� �5���NaZ�xvy��,�9G�t��a� 0��o���z��
 ��V�KO�����nN���p��1�ǁ��$�11Yf�0��k=~\���� ����G#	\}�M����b�)�YP�y6b���L|58�4�o���Ĺ!q� ��l���9 �V�pظ7+rB��~�X��A��au��M�~,���"֦�6̓u�>C+%n���uPe8ߜ*��8Fj�]$*�T���Xzkv@8M"kn'��μ��;��:���o����tv·g��1�7�����n�o�v�d�;���\*撙�:��fZߒ�)o4����3��6�w
���:9���TnA��A0������7����s_�G�Ϋz-���3����n�1;���<a���yd��g]s+x5`�'6��t�1�=�]Z�rN$�����1���#�:*m�h��:�2֭��f�m��k�N�1-?��1 f�2b�����c5�H�7�.{�z^����|�ߨC��)���p�25�������ܙ�AHh����2/��׹.�Ss7��Dn0>*���hO��3��e�>��քL��~�36�:ŞH�����O��"rlߑ�$I\P������3n�n��/˥�69�� U�{�{��슴c$���tᚏ׳a!�ٕ}�D�JM���y��!��k�jW�+&$ɴ��75㭇�o2��4�L�ɇ�)L�5c�i�	/����y��j�(%�A	�-������kM�;�W����۶�^��e��")�ݦ"t�(MBb�����5��WcLX�ȟ�����5��Ć�]���sU\&ϼ�X�Q�����E�I��O.?�|,'���������b����1Q�"���{��h��:�p�ݮ�ۀ����v���+�J3����C��1�n����N�w��:�,ĝ���wj��ct���v�}�6 *��-6������P�z )�Lb��ƻ;�#��Z(m�o���� �!�ފ�@;>��T�O!��#Bqw�xJ���������S:cw���^?�3��O��3z�|��{6�
��}ڂ��"�����.�%v��3Ѯ���-�����6�J��0��Ї%�b9�at�>�#E��i����e��sG�΃�Q�B��C��c�p�Ԝ	/и����~?�s���X��gSL�����q���/@��g��N>��s�%�%7�ae>y�wC]����\%�j��@U4"��軪E�:�}��_c���U�^�� �>y�Y���k��V��ۜ��!WI���X�3QtAE2�����j��
p���ޭM/*���D��$_@'d6!GB�# գ��J��B�ژ����&��T��ӤO�y�b�,���6,�D�X�uY��7Y�I�^|P .��v�o��q�Y��!�sSyJآ�V�вq�i����	��KZΠ$ Bs�Ce����m�ہ�,�'y��E�e����'ih\eEx������j͊i�1��k��TY`7��_�ܱDs'����k��)��3��Z���]�VX�$�������)V�,��2����3��2ޞO�[��N�f}FK�l�)�>��Zŧ{D.�dO�m���)���%��y4թ��np�����,M��RS(�2a6[�2{�Ӓ�t^�k�F?V �A�8O��9�|�:��W�[��$�g`�?o�LЮߤ���ň���U�?����K�hd��^�i0��ɤ,N꾢�K6+�x��'��K�ύ�bO����{@�E]�����![�H�1�x���o�w��#*R�"���x�|���U�͚�����G~=r|˽V�y���5�4z��ۧ�υ���:ևt�_��*xD5�c2��6es���Dhf֩�k{�t6R-nu����\�A� WfNܡ�!QS��i�Wd&��#���e?+aDi��i�8�=l-r��(�r��^ !����xa5%K|�b��d�����uW�����C���!y"�e<�<��c}���ü�"�n��|�K��a�O=��˅�}��+�q���ks�h��GSS����u2��NǴI�%
^:nF#�J$N���4��&R�ԋ��:�ys"�1Vc�/�}��H����V�J���g��N���P!x�������f�ݒ��@���+�7�F҆�K�ԆzS��(QZ�����օ����Δ�l徜���ApG���e�a�h|D���63IY]W��䕾��X�m�N����NB�N���PrbL��@��ȇݯ�GT�k��e/�&Z�L�j�W2}�A�a{�hk�ܐ"&WMɑ���FK�G�{�U��&CSR��4d4�K^�~>�C ��D�
F�i��/L���5!N�� ��yů�+W"�XU�p�T�Nn6��Q�*n\�K� 8֊�/Q2�8�s�ZF�i�z�#;S�&�]Ǵ1��I����1�NU\[��1����i�X�r�`����z[��sGb�;~��B�us&̐c�c	3����*Z2c�j!"3s��XZ�J��ae�)���*�PE�ᛪ��ײA[G�tu����-���h�Q�)�j:�̀yCK[�xxU������8��s���,���3mE��/�yPxb]��YE/����2)�_����;e�(+*��aB��o�����s���;ߕx�X���9t\�������G�-��a[.�K�B]
/Rw���|L�>zt�5��j��p��ɮ���p��j��~Sr.�B�L^�NS�-	-@g�t��L8���G(���K��^��KRм�-KMP�a� �*�>V�

�Ğ����"I�.A~��T�SMYt��M�U����;�����*f�	tLu��L��_�u­��-6���YV�"��X�P���A0��jkU��F#ZIU�p��H�^�P�Go_M���4�L�d#E��T����`5�^�X0A5z�d�������J�����6�t3KGm>�l�0u�l�YW���:Qa��\j��H?/^Di�8V�j�J�|�L�>��iĥ1�DL ;\'�5$2@�s����rD��ۃ}�1a:Ɓb��5��bs�i�)h�Hf�!�j�'j�Y��Wu�n~��O�k#�H2��\A�r(GMh	��:�3�͈+��,�>	�%�PZ� r}-��.��;�?����Z�B�\�
Nr�aN"��k��
�Ҷ�G��#��Ȁ��%-�#�Ԗ	�?�W¼����p����Vb7�3���<�ص����	�:��)��sczd������&l{g�釆�T �_�"��A�������el�c���/�ed�9I�2"9���T�:��4�I` �FI?{Xj%���ea`����K��������^0��.C�{�9����E���]z:a�h�Aۤ�	ݼX�$R&�!���y'�N\����PB+5��(��=�"x����ت{Θ�$��
�����z�B#�ōG�mY�u�^7J��B�Vΰ�\�y��G\�՜j_���3�S0�(��Z�]�g���o������W�D�{)�ѡ��`�[�T�0��n�A`u*�&J�s�p�v��2���ćy��ʐ�J���5�j@'64��y=�+���I�������Ю�\�u����c6�Wj�o{g��!��m�ɴ�R�����f$z�"���ck�����N�JO��;���RU��QǾ$K��׬�B ���A}��6�����i��h�q�H0�&�R�����	`�e6e��v�]0�	ۋ&�+�i��l���ٗZ!y�����9�t�ݼf�!!kvj�)Õ�h;B@f��Kz��C�\[�Kd[e�W.J&�Dϴ� ��^~[8�����&GI��n��W�cJ��
TB?��������u�����G�"p��^g���\O��/�=�K�9�w/W�5sW8=�#�'��I۲��Ns��V�q��w8�1���4�?�� 4s��l&5��N&D��o����n�Le���u#�g��V���)5
z�=�5({�~�w�R������s�sxl	X�߷��M��QA��y[Y������DKvX�
��F4�bj*>?�Va$��ܚ��� ��m%xS;��K�f,������&���/u dp�r�l���ײ��W7;{��7t��ϖ��^gs�W���r��1�}���!��*���^ë�e�Ֆl# �[/<[d������(��~x���md��UR}LQ����AT�π�uo�bm��]��oD�c-YY�(���`/�$4�lN�k�IXDBa��@D��w�RH��zM��
�"�Pm��4�[(�ӿ���m9�;*�����?�X��@�O� �'��8x2�3]C���"��QL�@[�<�*���7�l)g���7Ղ�Q!#��9gv�kHWN����iļ/,c0�����q}�`���&�`t2,ڣ4�y{Gs�����s)�f�f�!^�n��$�%�Gn�u�����+W���7Do^4�V�f8Fs@$�ȫ�4|d�l��G_)YV�gjl|��!JUV"8H�a�ڬ����R������B��[���D.���LW�?��Ҩk{�	\<���b��a�7�{�'*<��ŉ�(�u����"�X�I�������[�`�rq�˃��o��,���Y1YhZ���?�_@�~�p:���I�&�����DdXƽ�h�������%PK��\�hfҧ�|Ҟi��nM����co����z��]Q�<=w�Z\ �Q���WD�Eí�
�M�Q��c��Y���+��f��Hx�T�P�Z��Q���Iu�Ū���
�U �2é���7��T"k��o��r%-O�?=�� �Y �L�7�3bm���8�l�ԓS�&���,��\�T��%�x�sV����MlA�v�%n�����e�O�a�6�H�*��mG4�ΰ���U����p?V�w��\h����#��f:?8m����%ôy���Qw���g��-NX׳��|�;hR�y��.��jj�^���3�y��#��a���^�u��a�M���E��+���?����"��#{�ɳ'��mh_���e�� �S�����n�w�����) ��g͝�D�� >�cWo�n.y��s齃c���P�Wq6�]�ә��L�N�1.��zM|h�П6}K��O���*�/��r������F>��3�6�g�M/$>��[������0�j�Y-��p�3e�)��� ���2�B����>�@�E=��s ��𑯬���D�0�tF��g���de�x����:�~��&rOq:!�}��yuG.%-J���4$�?LG�v��f(SV��<#���M�ez����ֻ��'�G8�9�Gy��<ѩ��ɺ��w�7�^�i�﫴��,
��3百��ua��<�ٟD'r/Ӎ�f\��#Kb,ӧ�Y��]�� �6���~�\�8}�w�BmH�X�B�v���ly�Z��4U�r�LQ��(J*��D)M$)�=��i^:	0�f��4n��	ŷ�'
����c��#s���� L��j:�u#���I�c��-[�)M�+�	�S�7W��f�+�Ska ����O!8��6�l�����E�+Ŧ����<PB'��8B鲖��܀�(c��e\hdy>h]�	w[��8)�F�ƨʞah.YͦO)�B��g�H�G~ \���/������A���<���c�Q[f���#��0Ena�G�xz_�.Me�m�1��Sq���H�4?r��ݻk�l��Y� w��X�6�P�X{�*�<�:ND�ۥ\
��>s}X�ے�y�cNA[G_�>i=���,�f\��}R��	��>�|�A7t��ɣO~'��f�_�y;аew�˙�����X>�vή�kq>idMª$ ��%��N�TO�:}����`t�zʩID�sB��P� �{}f;�w>�{���*מ�o@��~�KEy�f����Z�_Յ��}�5��K�sfe��Jw��O��>�A���w2]RȂu�`��e�5	8��4��W��Q�c>0{^��q���&��A���S�}��5�}寍�]ڼ3�(�YY9�)�[~4؆?���u���� z�2��k8����I�~�6��]§~�au3|�Aq�אBq��H�@�ֵ���q�_��b��7�84"�, �݊~�l�"L�iJ_��{(j&N�(�k�5��oQ$�+,���Y�Z��L����Ɲ����V
]��#ۯ����7c�	������C�Z���`�KH�J���z⡘��H�L�GM��?�j:`r�uр�-$������g��D ���'��]���>A������v��'f×�{�nJ��b�)�a�[j<���K����n��#o�ֶ{�
q�r�Rp��"�I:h�_�����	�B��!�HkO�� �l�6���P˯������� �Q��$I��kYm��T �)��S�B2!G���\}��""�s�����/�Y[1�iz=w���*�ɓT#{��d�Ve[� ����JL���u˔ '��i?������Rh���f�D��װ��]T�	wz�,�/Bэ	���8�%S��p�m�����C])!�?�:4�0��[eq���N�/į*Ü}���٣�۶K�F��{o��Lؒ9��;�f�� H6��A�Q�KH� �"=A(�CI�]~B��v~�9��W�s�%� T����}���Ŏ8�w���F��Mr1��g�J�&G�a�p<����_���uL�f���0�q�Ň#��h��Gl���A+�4V.@� o �qS�gmㄴ}��귩�� ��A�0��5p��t��5uLȻ��w������ٞ�}J+SJC,!��9R*л��S�Yl\h�W5b�A�{�Sf!���n�y	 m��Cgr��M�5����|�u_*�
3�-J�i⥗{q3b��� b�_8�,�8�$e��5,On�.t�K��FT���c�!�O�+�-kV+P�lI��0M*�	_���������}q�5zWG�]�a�k8�~�� 0�q��[|y�E�(�m9��q�R�\<����\I����q�F������X��.�Qީ��t��d�^�ij��JSe�W�ŷ:/��5�_�}����M��k��Б���]�@�_��1֧��}�Z� .��<��*��eYݸ$�<>�n�w�&�����i�m��e�	�M4��|{���ES�!���������YÅ�N��#{�(�yiF(WbG�c������R��LE�3ң�"ٶ�k�阁�j��r�St�B�Z�<Z��}�v��L����އ|$�WHT����9�}����yԸ
8��Ijl
�u���$.����v����!���1�[�9&c��k93j�e:�+�����v!a�y���u>-p��D����Q=`yL��<�"QA��eRu6Z�� /���Z:����m?W���o'��%��;�GP�T4a�b��9S%k��(~W����y..2-_X#¾�l����1R�XgJ�|/��JܹU""��]F���E3y�'�u͊榫��� �����[�Bb-��CL�[�C�1V3�L`�����_�x/����2�Ê)�	�k@J�:�5)�N��#e;��s�!����g�����多�}�mH���Y���:ꊇ��m�F,��C,|�D�{�9E�7��up��G�Y��������t�m{2�-#�4H3�[ks��t�Ö�䳎�I\��{�:�z����ڥ1��uMΆ�OD����T�<�:c�{q�Al�Y�[kd�<�[�� A�KFH�Jn� &�J�>ANhվ�������r��oc}zJn=u{�m27aJ�b�:6���Ŵ�R��z�|��a^��^��W�RA>�%,�s��`v�6- �r�[��)���{;f�[�B�~�R��m��SK����A
< ZtA�b�.N᷻x�2a��b=���`�y�C(ēܱQ!���n$iҰ��Q�ءEtD��x.��17%$���썪P��m���rٌ��1l��l.F�@��#�ON���K?�o�)���_E�3��]�>1P��Np�26�s�#��RF� �J�
���O�3�g�t�\���%%g��3��*�^�����M��W��8��*)��Yԋ����,12�8�3��b�`%��p�R\��Ͻ=_�{�����ω6�{���|� ���T5�~_�\��x6*���+iq� ��2��Fv�N��%�/)���+�B>d�'.1�,�����.�a��c��\���1�,��U2�?��-x~R*������I������6���h��k�_�UQb/��v̼�ԁ�F̯�H8��ß�9��㉣�
5����l
5M���ӒM�w$8s��A�+�u�X��*�k�NH�67���=�*�������kԻ�V�u"_��qV;�~6І)�<�Ȟ�lj���~����N�6�A�Ϭ�݃����c��8�HB%����;.��%[o|w�{7,��#��L�ҕ%��/х �ld���3]}aT#NC��j^�3d�*t��ypP�\���Y�Lऍ�K�x�h�~;��1�(�_�X�1��쪼���ř���;�0t�W������^���I�ܡ/e��9<ѲXdQ�$���\IG��D΢���ݰK��`�@U-V�b�dH�"(䟒�͊z0o�J�Qe�J�u�#0��v�4�%���S>�í�7�N�#�K���
�ڝ���h;Vm02���Y��tJYH�z��FD,��^<���*��m&�]++u�a���;4=sV�hN~ ��Y-�[ m��;Y���f-qV<:��������� 0�s�����h:{9qz��fGy�>y�����5�I7� x�aґ'�K���X* <�&�bl�(�u! ��C0��hc�U�����|^�G��)�v��΃������UjO���'|�4��_;���=�������ņ�����\���y�O6F/k�RTiKQ�a	@�P��/�#�?�*	�h�q; ��C�q��S�io� �o�'�J����^��l�+GRrn�y2�V�#g	eN���\��;�
x���߄M�t�/<�D~Y�:�/F��כ]{ϚUV.�
/��E@R��k���-�/�u�܊g�ؾ�x9�`��pF��O�t7}�)�t��hz��΍�i�XE��k�
4��X��K�;��Ʀl���E��B���E�h��~�T)(�(S?�C��2OPO�E��v't�g���sg����a�S��ї��A
����X~/vhF`p�ΞT`Q1�2U��!��F��3h* \S���{��i1���Ն�e-����v���L9�fI:�yIK�dk�zo�<������?�\��{����#�uXB+�!�g	>7�m�&#��PY;e�yPƞ�jӨ8�ek1���p>�=�B��"��3E �J�U�(��J��9���_���g 9[c0n����i��ۼ#��|�"����.���"���7�ö����U���Q\��U�����x��@U����hd���r�%�l��~��0��Ҝ l14���xT�w9K�� ��QGg�j�vLjΉ��ߤ6ْ�zS6F_-��`����\wX�W�Z<~���x,-L�:��,�<Cr��ҥ���,�_㳗=eɞ hWFN^��2�2�
~vK�J"<��hl~�)_͆�D�!����f"�C;��P����V����zW��˾:�J�x�G�2.3�'hg��޴qF@��#����Ј�����}Mt-�'`�S�S��@;��>��O����Ni�8��:Z�
apD��u?�Y�N�!�V@��X�y�S9P,O�u��IV�	�'Oh���Z�k�AeZt�⹈W�3��l��O��0�Gm��WOf��\� ś��4�L�!6���P�0b���X�8N�ڧ�{Jx[�gi�d�q�)�sD`-�(��XR���w��鼉ι���H|��x�T���g�yY��k/I`�A<ξL�� ��_���\��O���Tsd���@h%�a듗�/�!��O3J�G��h�� ��p:�����NX�\Ãn�?{��>�l��װ�_J���g?<������]����آM�7�#�����H# �|�>�Qv�ٿ ��Es����^Wg7 ��Y�\����Qwʹ;�W*g��?�c��M/�/��&e�o�A��ލn�?���ɨQ޸H8q��x�$����ho<�4�d�1G���hGD��_E������-��Z��Lwe@k*@Y�R�&�2 ���x�^i���y���e�DfZ�W�q8Ҝ���5�����\���j;	�Tg���]�%��c�cZ��^d�9�U�Ԩ��i��$d���N�Iy7�ƖjI�̴Pl��	��a��g<���
��di�E�8�$�<N�B(s���>Y����To�r/@yY�
�r@�!ن���P״��a��3�0z`;����|͉FH���V��xY��@H���L÷0:>�f�
�A0�� 9n��q>��5�
ݾ���ޅ:-QC�������G�R�_P��?�`#�G�$�~���}!�+Fn��ڒ�+@���:f��Y�p	�������i��D5���&ް�3V����^�vPL��L��4��3_���CYְ6�I���h%��y�W���;��I!�F���6L��� �Up�7��8�������}�����s���f�Pa��D��E�H~ӹ�ko=SC>���jad-֝�X�l�Y,���E�\Af�[��l_[^���;l����ckVg�Tq5����9�I���5k���Q��k���$}ňPk���Ƣ	f3� ��h�Ԝ"�E�,^Ҟ���q���k�!��h
�,
��VH4t�-7)����A�mC�b^E
Ҡk�'�V�De�x=h�M�չ@�52�V�i�ݭk��A����>�U��P���e��{�%I���AU��3�� 	"ձ���Hl�_i�\(OëVRPJE_�-��[��XS�Լ����zY@���]�t��V>�9����T922�^�v�0G���֏��-�����nL(���X㴱Rzl���2����d���Xޔ��$�w�B�HG�����ݧu�p���;ĺMr�٪���q|E�d��ˊ�A�r�y�)��g�N�����.�i=`����YC�o8�W�z���-�3|�i����و�+Ti�b
x-1��"N�Ges&��6o��}�9���}AI�3���c�u�%�ؘ�k4ǳ��ۯ�J�#�m羺4|�4�2�"dd�j��D�����Zn���j�le*
�r�:[y��Sa~�T�'�k��s0��O��O��q%3�TW�f��{�w��u�9xe@����oyj��4t=JUa/W���gy�aL`�|�mЕi	��H�>���:�����j!��<aE���f�M��t��H�z��p���/0�	�۬w4.v��q4|s�,EE�z�֏m��QU$���[�R�5VJ��]����D2C�ZX��42EC����Mxk�#� ��%y�Vr��������c0���?�E�cɤo��D����S����1N�lϥ��(��N��c�����ت��������6�� ��%~�v=u%K��'�|���±|���f�t
�jv�gv>c�P���p%Ń*B	x�@�Y������˨�a�(�q_�2�<�߅��!��H�)���
yV���*�,��a�T�ÊM�O'�`XƵ5!-?�� �i�s1]ɇV���l�Pfi���!X�I_�چ x�a�R(&�؃�U��y�4����I���Ϣ�t���V�N���n��&F�J��G���᷃������T�t��5�����m�۫����a����gV�a�\uaB�43�cm��T��|o~�G;�/�����it0x���?��3Q��^�ϟ-�p���a�*�����W�k��5�����cVW�7t׾#HH�Ub�JHkO(��xH�͎ 'B�̲k��e�nf�������}�0Yo8��E�yӬ�1/�����ئ��s��]�JK*�y��$��.��J0�����P�J7X�N?*�����u�yky��J��I�v˦l(������l#s� �ȇ){{"?h28�S�	�(ۭ�|_jP.�<�������K&!Pc��1����L��Fn[���tZ��c��7졼�n��y��U@��U�����/�ЌI�8��̿v�]VW�y�\Ri'�
�=9&�J
���I���h��(f��|L��v|�倞xr�{^Z���t�����)��q�D:,���b�W�2�!ʴ�?�5D��%��7�u�IJ�*}��M���=�ߥK�x>C��Kꈉ�I�xn�N���{��e�LfpϺ�ț��WL��o9��csZT�������T?X����𲶰�I�[0\"���0��4�[��?�{L������^h;3�y��#�eq�������p�+p4=�� ���<��M��щ�o���2�����x��5�r������mc6{{�o��pOՉ��s�S��D���wxē���m�J��=�� ����D��檨�hDq�{$�$g �]U.�tEs�恆Z8�׋g9r�߸��mS(�&�qC���T�����W���u�F��e��q	*����,��Hg�Ⱥ�/�:�������RA�U�?�=���O�B�$P���|J��W��ʣ��3ZM<����$&M����*�D��
���s0Y���5!���_NO��������Y�U(Y��s�f��G�V����m��WW̏��8"_��w�yNs)�c�g�I�3gO���6��i�E"��� �v�oh)2S4���l�yv��7|O`�x$V-)�KR6b�u���Z���|�O;'x��/�_Q:Y:
c� f������0�=�ݴ����3���wޙ>��v����C���7B��P�-�7T�����^�`�i.~��]�
�)��n5���.L��˭�x���(�Tp��V�zG�g��NT0���;Go��n��V��S�\]�AM��X,͂����È`���_��Z6cR��^���8wpM����˛z_��;_R�7��pQ����ʋr�۷�&W����? Ov8�[a|�w�{d���x�7������1�P�>���m �8�
V�R�/��2J&�s��A�ѷ�����Բ�����x��>��B�e�꿆�A#�u�5L�ZJ��x�M�j�P� t������: ���c��]�
x�L)p��r�H8(�5��{Au�#_�4f��W�צ����&L����a발� �l���rk��4h��ׇ�i��,���=^^�JU8�ګ4��ӏ�8 5J����6���a i3�ԞT<�qe���.I�Wb����ҧ����8�0��	:���9����=��G(�4R�?{0����Z~���H�c; ��)�sY[�|(�Ą�zI$��ݰTx�A��]��[x�����%��z�rֱ/N$S�����fd��
�-x����ģ�zt��1J�� �n��p�#�m�bf��o*��p�?�m�<<�$&6T⁀��AU����Sh��/4i���n8S��K�~&/hm��twk�Ԭ�e�0���SRDk��YW���P��&����֜2j|a!�O8i0��s�S��.0G֛�p�v5���=�ƑwRw��}k/��h�]�K]�/~ˊ� �E��#?ʅ���������0�_u>U	F��P�@�f����U���/K=�I�>��
%��y]�wJ���j�?�����K���.����D�?k��!��|BC��6F�\o(�\v�a3�Ǌ69����s�
8��Z��ש���.����y�c'����	c�t��G�bԘ�%�6;_�^5!�+M�2�lc±��"'�%�<IQ�0 �F����d��N�H�e�IL/9�G���,�����Y�]�����ٍ�fQ�X8����o�n�����@�
05�܇�)`�S���k��+�_�+IU�[]���s�<��Q�r��Q��-G����VH��� �d�K(BA�ͨ����c��VZ[';��Yp�zc��d�7�M,��n��&��qD�iţ�����I�}%L���_�>���E-\;��Jg��c>��iQ���.3O]�>!���F��
vh-( h����� Zb�E�em�Z���zd|Gi��h���N�C�"梍�B���jr
�<xW�^N��[�2}��ʔ�a�{�P�Zp$�U���K7�S��Z+3=�p�)O͗�=i��/��:���q���7�BR��͖�N���~���}������ES0�����჈�)��d��
i���Q��{�
�!|X_�j	��$y|����Rk��pȻ��gE��4��l�'��My���!�M�}��ʅF�2�@F��iZ�r&����
7�X���@�R�Dg�l'��&�9�ƚdʋ�c�Ш-(���Q�tR�R.�I탄���e[xD���(���������-C�V�tb��������ۈ�d�p���Jb_l{ʼ�Ƞ����VM!H�R���p��?�3��c&e��6���o��������\�  ޲�Z��'g�[��&/ՙ&�a�U�*id}Z�u�/��R�h��"j�M�N\���)?�t���D���z�y=B�=����ϲ.
\WR���9���Z��;�4[W�EctWڗE�r`X���]��ᣲ9,>6X��,iq�Fu)3����%�睇�%{O��[��}p¼=:9��ߡْ≗�z< ;鷡�X�"��+_�꧁)��ᐣ��cv1��-FT���������l��2
�
����!ת�^mz�2�̾Q�,����'�$�6=o�����ʈ�-��S���f��t��@��߳)
I�:0"�q�������u֋�G�l[��O��T::�|���[P���'2*�E�(�_YƎ�_��<S�(ۈ�PĚY�T���o������!��C�e5�Чh�y�8�d_�����}�@�_������+��\������I_
�=�PR�p�J$ 2Aw�r�u/����Miy9n��I"t,�Y�k��.C=	�5�S�j��$���>�s[Z%{�C��YͯN�
�F�D>7k�v�=�"��D�|å�����)#���h
;�x��~�?��kf�щR�n�!5��X"C�����!�.-x���l
;��]*f^
Ɠ� ��ERA��5��Ţо7\l�_®i��l�5�`T:o�D�Iŉ��#�wޭI�������3l�,&��tq�$y�0�o�*��xk4]6��[�����p�%���>3)JqM-��@��q���2V�*MY�����K��8�8a`w���1(8Sq�I�~4LV�>3ys���S�؏���E�< ��!��N�=}���'M}=���П]�<��A+Q���O.����L�n���ȼ � [�H��Q]h_�"��{��\N�0R��S�ͽm9Bg�%�E�t�+q�/��k�(}QM{��+p���P�=nƶ�M�VNF<��W�%���A(�[�u��3i���F]��O�ʇā���d�X�9Ol���y�F�m �~��5���u�`�G�:�`.��!-�9,l�Ԓ�Y�!�򟓥��FQ�����|}<��j(�ɕ�z�K�8�Zn\Eb�!դ�~���$S��n` ��kX�^�d�ZGU���D��p��7_M�b��5XֵU���͹h�1N������ �5tX���Li���!��Bo��9ɆC����I��&���UC.=�Dǃ?�wwxCby��U˶]���+��$c��1������x���
��-�]����S�#�눪bFx�XŒYﺼ���h�.�n�?2���ՔOlt4�Q���q��Y�/�����@P�@'0�l�u	�.�$t�a�W��U}�Iox�}����pyק�+!��fC���3/�Wl��=�g�����|�W������NOl�f�"��RL�2݅�Y�B���A��xO�ɬ�EM���g@�R��[L��2�fe]�֤Mά�hӠ��UjKfr$'�	��B�l���I�#:�np(��/0�'Hl()�1�xb�[۝DI؂�2Fݏf���qz��ˑM�"M`�}H�X�8�9��>q�W�X�)JN� s�Tu�g�{��e"�3�;��No$����������K;,�?pL2�eQ��g��/�(:o0��`�Ƀ)�B̌r	���%���N鮺�P�X�vρ4C��" ]�o��cB��
=�5���<��"������t���� %�9��1�?���v��BA�cI�t�S���s}�O�y�w(bi�)���{����Ǽ���d��8����b������3Kn��>m0�t��#z����K�o�����YPgv�q�n6+*����R���Q��2�]�&Ħ}܍�#��r@������¾P�H%EPz-�d����=|�d|j��c23��m<i�Q��%)[�Io�8��*<X��E��N����{��s��S�B���7O��x����h1X����q���>������z�w�B�;�W�.E���W�	+���������<Mv�7�K-a]6��{p�t5����Q�=39����q�ן�<����\֋��>.�m@�H{ �o�n�(�|���R�/l��B8��R9I�ko��˼��J+9�#����5��{�Xm�4��e/��n9�*w<����[���@�s�0zu`�����*�;=8�y��1�}|*3hi��]c���`"���]Ά<\�O�e�����S�уgA�#�ce
��y��	�
�6�"a����2~Lb W�ĔZX�=t����۸YI� �S�g��l;e�3�D	�)ϷU9jB�Ur�������v �W���2��~''�V���5p�3��ö|:�S�vU �ܝ&w��g'�ˮKqcK���V$;R(��7EH_�e�G�a�t0	�"ߏ���!1�q�)܄y���a��j��	�*��,A.|"��0�.h�ҭ�����tF�N�u�	���K$����(���6V�0�������=�,��0$B3 5��8�nhƿ���G1'�m=*܈�'��)4��`]^�VF�O���!����Z�dD^2I�݂�|��lB���Z!��[ b���1��\ ��1��`��8�1[ob=�6eW[Ͳ�B�+�0�)I���d����|n��(ظ,,5~M]PK���ҧCm~�S�J���z���v(a$�L:϶�3,{Y��x���N.	m{�+�����3P��(�iTx���8%bm)�w���r�N�[~+��O3pzo-.���s#�(�g�X�`�C��[���V��d��2�ؾ��![�6GˊUbJ
����'c5�l,D��]2�t7Q��}���јD��	�a]���4�Q��c�K7U{s�h��@���Tu|$z�e�~Y�0�T�?n�C�r���\gm�1.�@��-o�j'� �a|�	�p���K�E�ͩ�*/y�9#���C���"�IN�GM6�v(�
0j,���.�m�n�(>Ĵ1�L�ϱ4/E�p����}Ʌ6\��S^e����TD�k�gg��O�	�z�%l)��d#T�nRG�ɏ ��zz��Ѻ����ު@�>P}W�k�:�����%ҝ��y�'�H�vi�l2�j>�X	ʺ�pjz�F7��5���{���HO�K���3�u$�
+n���n�8�܄(����UOj�q��l���w�S$@[��<G�)�3�������]};j�j�H��I�Xs�i���9�*��1�qY���AC4�YI�d��8�bA���4$��XD�j=��q�GH'f���>q���}󈍈Re���ڹ�hT7� /=��+�"�q]��$��5 ^ܿ���A�i��bLD�x��(����OX��x{�r;蛴�s�ǵ��[#�7A�v*�@�H��w>��%�`�H<�r��d��Z̼v�n��Mp��_�B�+Jޟ4��J�U�Y��tr9����D@e�=����艟33�B7J&Yn��^X!����.�/饐k��uI����m%/�s�Ew��[iX���d(��uWy�<o�+�1�t��C	�\���c�~�d�/��Ǉd�l����bI�`�ԙ	��8v
��M]U�5]���YO��0�ٗo_��:���&�~�s��(UX������=�l��f�<���-X�\B�,M��� ����K�`Q���܋_�N��9���!��NpSx���Q���@R�\?R\Rʰq<t2�H���:9�Ayyq�"��#,&�?I�Q9��Pb��=����ᠳ%I� F"M<+;G���:*�R�`n��isS����`�-�	���Vn�L�T�O!��]H.e
��-1E��k��Hܨ�_(�ǻ8�_���g.�5B���y��<��U ݺ��L<�\9T������Y����ʛstd񺕓5��Uh\`cCT6�,�bؽ��9�HÊ����4Ͷ0Z���]�Z�,�{d�8k0E\.jV��-? 1�`e�0�eĦ���5�����<�0�x�'��NA��rhg1��S���]R`n��9�%N�Tq륚��L��4���=�����|ӌM��#���Ww?�q��=f���-��|��N8��H=�LT8A��o;�i�<0��������S |�604��ʆ���
X�y��FX��M�K��x���x̱�7�j�k9�B�ciGZa}5̥�V�]�=��g����ʦ���d�b�n�n[�Y��M�<��AqYu����x�J>�GI!�����C�۸���0w��wY�M�
ۃ����r/� �d_�J�#��h�x�?F�V����V�#���p�p;��n�ww��1�Ξ���68.���Q�"\��% �o�\	�@c����J�1V��߄G�1st8�l�*����S�������O��p'D�a<��mM��f(OJ���}��G�&Uj/���g��y�N��b>P����p(���-8Z�+�@���7H�.du����ږO;T�� �
bڒ���N ��L'�S�g�ߎg�Q����-o��3�.�d:����{����|�!�aU�3}��0dmN�D����݇�1�����%$�Y���Kn��dv�B���v��en��,Ck9$�6��џ$6e9�����~̳�y�A����\g=b��3�X��ee�qBT(s�M�DS���](q�ǱM�`��&}Q���t5p�<ڊ���	��;,rl�VERh�vܴ��vGnY;�"�j� ��j�(�A�?'$|c�����u|��*��U�m��K���\O��}E�y�S<Y8"�vςJ�U��:�>�8�h�/,' gZ���vN}������&�X1>hè���� [�&0�\5��=��	>��4�*���	��RO�R����7���_ه�J 4��@�p�v����-���%�Ǉw,�U����+��J�.��{K��vJ6���'. %>"�+f��ڏ�8ͫ�!V���W)�Xw�]Y��H[��<��uWe��`A�W(��6�7d-�\��Ɋ���%���}�y9T��r�1Fqd)X$@�U�)���<��~�@v�}�Rq��� �.��s�D����놃��[�t��Ս�PɅ���fyR��|��(�:;�iyUe�e�!���V�l���+�����3�a��2"Ĵ��Jʞ������㪗?.�C�3"�n���+����������U�\
i(�������ׇ�����j�	!����F����׸� �v-v�!䂸7��e����Z�&�,���%�ݙᶲ���Zf��pB���ˋ�Fͺ���m�\a��B���O�m��n��}'��M2����M)��Σ���_��q��fp>��2�݊\ ����W�#d)��I���V&j�_9�$��c0>.��U^�we��V�u!@�2��x=�h-�����pd��x ���k��̐��BX���D��"��(Z%��T�fW�L�'rF�j��p�@7H܋q�x��c~m��1w���?>UQ$�f�=@MD�B���ot�J�G�${�O
��J�cTL���#[w�ǔ��ZCe�����O�xiɷ��ͤ3��|}�1��V�T�Q_	�����J#���!�����k�FD�m��NhI�{H>��.Y?���aQ�n��z��o+u(r_!�!>�_�8�#�G��� R����
�ҷL=�W���L`M�;��fE��ňJ�4�
��tؘ�V��£�NN$�*����(��? �m,{��uv���16����qCH)շ&y�U�1T��H���E�_��� ��>!��b���ϿjCo����v�*ǃ���_�]��#<�K� �&���,c�ly�ڕ���\"X ���J ����'�n�q��"o��Q-���F��V'�s;�d �6��:@ iJ��2���7�%�3�q�Edn��F��C��9��8��$��M�͟}���l݈��oNo�lu��e�2ƻ�]5�ɎO+.\�ш[�5�kqi�d����Õ4 ݷ��^ k�"�Zm��������ϫ$}upo�j�vVǀ򰫨��HE��(B�NTO6.�C�q�G��6
S)&s�X����5&@�2�lZ���֌���1O$���k���M�`�/)S�Ԓ�~�;����rseLԈ<�">rVM5�)҅Y�`~��'N�dR��f�����1y�O^��Hj8�}YZݫ��.}Y��@���j�^3RC7�KTc>	���vb}�>�ܙ��S�]n_wP
�9)���P�n��Ƨ6i`��y�$�k-~���R��NG'.����j���~i�A�%����}_�n5sR�-��p]T��/��z�Q������e��9w�D\a��;̞nh�7�[��U�A>WK�oɛ����"3�Snr���W��K���ߙ�;!�1lB���=M��l��Q�,�\�]g�3�vB.��dd������8v[%-�4�Xi����Q�y��Ѝt����'Vǣ�ѭ�XvE��
|� ��3�^C����^��L!����G�)I.i'%�5�_1�#'}�������Gh=%tSß�`��Ud�S�6swm/��Ng.q�+�7`&�#z�4wn�����R3���6X�'�{6��_�3��q %(���.���\�|>�EM׭�Nݖil���� ��A]�0����z�
�ߗ�:yMU��/썳�r/�]�g��a��c�J`xT· H&Cfg?�jcT���'R$hxG�_��We�u\�p��Vk���(��5\��%��։4�PU@>B��������Y������Hr �a�as���?����g_8'�Ѵ���ivI�#hx���c�ȸP��H#l�Q�j�۝����@�2q�5�hk�*��D�G�K�@:���M�����ZC�O������88�L��H�4D["�	�i˨�4�����s��8y>Qߪp!�ڎ����5C�2�xKM�(3p/>��Q��}��+�e�ˁ��̂1VCaS����L�v�R/���BT#��W<A�*�ٲ���;gI��	��v-�=�.������_W7��ఫg*�;��j�l�KJ��^,(`������fX��V�Q8Lh=��4�ݚ����%d��@mw���d�ָ��FO,C#-'��_�𑝸��('c�dɯ����k��i�-�I��a���T3?�J��c	IG�"mX��V����H�(.���MJ���PC�<h9�ꇘ�;������e�������T�����i����Gˀ�h��!�\/�\0E� ���pV撼~(Z��)�Ư����Vt<��c�5��	��)9��|o���> ��lW����x�Ê	A������y&
�J���ɟq澼c#jojc��uJa[��v�M��~)� !�]�P�6�۷�x�ь�6q��	6|�
g�m�+c+X~��d:��a b��vN��:�cI)���b�������9�sN�ylS@�2'�}�����R�wl7���bc�p��"��GUM�`C��m3�]�V����w�yN�]��4����¾X�~pT�G�q��a��,�Щ1�%��T�@Q�9���S��e�2��;���� #���<�͆JR-z��\H��-�o��<�''Sj/�����E� �e�ˀ!QB��nd]����dm��Jg��%�|��H��:��j�#5�����о��qɇ�'������ꜝpx��w�]��Q&��+I����bw˺O$��.8۾`�me{Ӻ��@BԌ����oL�N�� ����L~0�=�)x����*�%��'�M1}`���96�~7*#6���X"~��7e7��/F�g�]Lͨ��P�D����,%H��ㅏ5�3�/�ǖ�����au^�і�̒����Դ�7��&;�츣��s����G@��Cv�Ƅ¨���I&�Mõ�}�����R:l �q(�d�� lD
��@R���:� �+Q`��k�׋tV��X��s�EeZ~h��mZ<Ƣi�G~�@JB�""��ӗ�&�T�E�����T�u3q�q���C�w�;:#/����9T��F�\�v�{[}8�Ȼ0���e��-`�U+{�Bf�X]�2��ע>�Q��kG��+����&̑���^g��_҃��ԻKk>�x�d��,��Ԏ Ҋ˶���yeY�G��D�#�y������ғQ�����g��:$螾��m�H&<uqr�lkA7���H����c��	�Q0r�&���(����Lo���5c@3���"�j�@/e���H��o�$�,�l�� �����)_�-��AS���M�fV�9�����1Pρ*��c�Z|�����H�\�~B��hm�L#����C|��Ir����h�Q��<]r�_S���1��NhuR�T���6C�65�����[��ge���$�@�~�`��(x�}Z�S:�*��BD���2�Z�cL�
�%`/�!U[�eM:ء�F��yR�e� �+��锠��l�z�����a�*�;�*�YxK�p�);^�
P"=�>T�����<V�.���q0?��5���e�>V`�����ioJ0�g���1��"l�d��xe��Y�*%�+�b��h����-N�5ݝ���h���0��Y�p�-IW�����3uR��ѥ��*0���DU�=&�XaH�#c�mϡK8�󋝵2(�9�ԧ���k⢝����i]��S����P~�E?�^B������Eέ!�7A'�a6|p;�_8݊9]_jh���4yF�O��:� �Z�\�ِɺ��.a����礐!�Aqx$���0��|Y:�U�r)��o���cI���Ws��-�0-�jH�T���E��r�b�F ��3r�Ä3����^�8����ztRi�-.��CQ ö����I]?�w�w�и��ɑR\qro."��b~Q�s;��M����q��$�W�~!(`%^#w��sd��*-h�_��������X�8��,MU[�T�H���������5�~K��n�W��Ж.SJ�s!��D�&<�����Ş�^��no�P@�� �� =�E'���	gha;�� ]���_^eڋH�|��,^��Q�8PX�$7����_��3@��~u!Q1���:��m�p���ө�M[��0gf�t_��p����}�XL�t��r�����Z")=�E�"3��@c�#���P�`�T��R�x�ș�����e��qN$�<����m�&+/#��V�^dN`&��v�*���T�F���EFL���q�ݧ��1�7��?�LhMf;lm��P'd�3c�G�8|Xn�)t±ޫ:���>����&��IF���e��������x��EQ|�'[��>;�C�r��)f��M6��� i��������@n;�3��yS�⓻:��J6���7s6���jÔ(���
$2�@*{���p!1�CVm9:����p}zR믝�{N����m�	 ���9w����H��TA}EU ���刡�Oqgd���E���f3\Qﬧ���}8?Tb�Mn{�T����mof�U�<s�"y7LWn�@��P�P�6�F��ml��.���<G�j<o��?*������>E�m=AYU��$�'���&�W ��!��_��i9�]�.}R�u���Z���?7���M��`�-�����`��D�ǁ*��]5�C��n�V�L�9�N���"@+�C�]���t֪�uЪ
b�a�B�3�%'ר�h5Չ\����cj̯n��dk61"֚}�%�.&�e���[?� g�su��Y�{�퐞�V�W�!h9��l�@�8�o���� ]��Xˑ
E��������JK���s�VN���=�8���5ȵQ�8,W@_�������uf5'��J� �d4�s_d]-y_��<�<�ç�|"*���j�D�Xi�8����ĚyL�/�Ye��F&W����'q���f]L3�<V
P�Fz�����JE��Q���l�|)�쭮�b�\��ҝ�Ҋ��r(Ӱ���r*���>�}iij��>�X�Lp�����e��$YR>B�!�ln�	��Z�WK��ܖ,P&f;���z����-�?�ιC�V�X��k�p�C���UO*��+����2&\"��
ݓ�J���Qa�S����\��~�߼���C�&�*�+/Dy<4��<��VJ��O��;T�8sN�v��u��[H��^9��2��
�k�'�ws0���S��"-�5Sk�vΑ>����{iFKu�MԒ��L%��Mv�!E�w梫��4��Z�٦��EG4=���G	Vb��kО��?����{�$l��.���8V��."9H+c�x*�pSuk�q����2�qTj� ��y5ȣѺ�'����b���D��F/1>ކ�����*6��f��L�s�H��o�����+� x}J��q���A��(���]�s{zyug�H�Y���#��3ZS�,��vm�>���$��������5��q;����,�T��L�Z����4S1�G����\���0�Ng��=7,�7(��R�>��u�褦�CTք�����Ӥ�k�(�Q�\9��k�?����
�m�N!%�Cwj�	�V��%J�vV�XRc��������g|���!�ᅤUl�1����ӧo���`q�l4OA�I�W�)���I��6�q�\r a�Tf��Ui�)�
ΙF;o�ٙ���p_q���X�/�T{�<1K�1{O:�����\��g+�P�)`��I[�q(b�gKR.9ͷ��F�W�e�w���E��pk�&$��z�����ӹy��~ �cK�X�P�w���_g��Yڜ�"�-~��s�αB����j��x�����Կ��F�����w�]嶿۸?`�?9 ���yj�T_��a�Ƶ��5����!�ʇIHo�p�c�_��rM��1��sw�f0������oE���ʤA6$��#S�Ú����8��4�~a
R�e�V0�8z�w}�8�jZl���'��Ys�R��Ά`+\R�Vo��������H:A�"�i;�CETդ�	_�U'�[;�%�B�,�lcvh2[5���+Q�މ�/C�ֿJҿ��>Sj�ڳR�g[b?�W�ه*Z'o�����ڬ�@*jN9��t�U����~�Y8^���cN`)a��)`��`0	���Sr������
��+�Z���
�O����^�"=�A�'Uz#�n�+�رXa��pRn�W�f�C
�*�7(Q �cF��
9�����nڻ��$�L�Ue{m��.�`�9�QP���&����B3�ö�]o"��_�J����ieg��F�	��/"/Hz���)#�yxݱA�h�U�����u�)�ɍ2w��G��!�[��Ŵ�Y=>��)�6��e��V�:�6
���>7�`p���+���>�k�
��F�U�l/���ASh�Ʊ�f�~������ή,E�_���V�6�y"9|��*���=�cխ�D��0�.�H��GJ+g�p�HD��@j� ���,hsh�gݯ[,3��r�3T����m7~ܘN��}��T�⍼��Xt�\ä��P�>�����*����t*Z��g&}�du�0u�I��k� �v�� �*7��~�c�l\�)���U��,>9����"�u8�x\1v�p��������'5�� ؞�f@��Z�yH����;JϤ�1�͜����6�A�d��r채To�z�s�#�<|����5��[�S��ZP�'�o 
�D�7�~a+dy\]�1�9�BD�'�o^1�z�p=��&�.-,ˏ��h'�q��cl�>%��p9 9^���F�Ҷ9��8��%��<6\K�������	z�`�o��cN��'�Jˌ�;՜�t-b�ƸY�,)S���<'��p&�+TM]
%GW��<��+'vPW|m9�7�kYGnf#������q���f﷾�c�9�	s�SG骤f�=�o��eNn4K%���v�M�6�j���h��6<U�tit�P�,=I���ڥ��,�J܃���*�z�iB
Em$��nv���ct
:)��W�E�n�Ø͉��r�9ӑ���ְ���4�i�>�yѮߣ`�5��U�}�*�2���ϖ�kԃրyhOH8���Q�$��r҅�g�>��?�\I������Y�J����M߲��0&[s�H¡-�B��c�|�38B��i�����8�����º�sbU�A�>����卌ɿ�e>`�ۚN�ṳ � Z�FƔbQ8�0���k�ps>��o�2�PB�^�&Y'��T.خ�|�:��5��[�we	o�G�;/L�v�WY��Q"��xڟ�Zu=������̈́	"
f���.������y&�%گ��d11;Ec�LН�����Y|�F�Rȅ�����׭�"�c#�F��CBAH�7�o��ɸqp�D�%� �z7��q��uwL0�%�NHw�(��1 �rG��<�Z����b�4'�-�[�c"�3J̊�w^�<k�۲|�W˳4Ì[U��,� R(��P(E�x����;2��a̦�Z2�5$�%�|���`�:��܈���>��/��XLh�^Hs[���y?Ѥ�k"���+ŵ�ƻ��2p�L(	ݏu�s�/��i�x'�����T0��a�WO%���z���ʯ=h�Ӊ ��[X�أ�gW� ��R��4��FB�k�ù�����E3I���Z���j�Z��T�̉�߫+�Ƚ����1��xyA�N$��EL`�3�6�*����%���a燓�B$1�����7���0r.V7���i��\B?�.5�[x)[���=����R(�r�`�N�z�Vk9A�t�Rf�>
�i���j)�B^d��N*t>WW��l_��zD�i���@%���x�9�VE2u�9�a��m r�Q�܍���w��U��6��>���k��B��OZ��&ԏ�d�5���M��z[�D�O��q��������K��K�s���N�DY�U�m-�|^���Qbh%i��ƚ��>"��1s��kVo���?7m�g�����X�%+5��{Bm�nH��zcφ�N�	*��3L�NK��>��O��K�������@�m�Nz��$"4x�g_��,�p�'5(RA��6���Lx�ͼ1����U���OF�N���,�u��w�
w�]��{��J�k����wc���!�8Rm:(�g��'-��4���Y	[�"�x�3�{/�H`�ӑx���H��-W�Tf�:y����_�!�Z.���ȡ��o�Gʀq����ϝϔ��4�o�6���tm�m�C��ţ`�#� ��T��y]»RmO�W*{��̗�|���I���%�f��G3c�hO	��F��?�S(�M���-]���S�#[
�C�z{�7�i'�2�4�Q=�CNL�}�J>��L��HEM$�*�)�Y���M�bQ����x��H��nn!���5h͏Vf����&�d��?��$��S�d�{���V��c��=ⲩ�7���j��8�?�(֓��I=�ګ��yψl�O��Me� �4"� ̶!�V�t���ު㒂v�^"GR]���D]c�ɳ�0Q����ΤBg�p��!��,���|ق?���،-)���Bb^�z�v���>�d1�U_&������7��-�&g�
��v���iLߓ�V��	k�n��؅C���ۢbS�9�HR��x���x���>�:EmHK��9�cZ5��o���3�oن����#�<U�R6�-L���%�~\�D������8����1�4�4U�+�C�f�hx�~����gH���u\Gw��ƘG6R��MV�� �S(-��1N�S$��St�;��q�5\��d`h�I�H�JV�Ȩ���jV��d��0�Ρ�7<<���'���Pe�șӖi�A��6���,;3�R��0���M��(3Ayϱj�G��J�!�fjR2��,h+6�3�����U9��JJq���C+�\��%�Du��e�D�T������U{���I��/5���^���_-SL.������t�g��.����?TG��;C<����i�J�p�e�&T�-;m%.G�~q!��n=�z9:�?��C��Yk�\�lT2�z��>�74*す�X�O6�ٹHߟ�v['PH��A�Ra}�6yM2�	�M�^͕[����d�1�N/�z��srp�Ơ�Ų�5ٗb�m�I�<���f�eWۨ��D��������߹���մj���~l& ��4}���ݝ�J[�I�|��9��}29�Dc\ǥ�bN������$�[w��n�^�N�h=EL3�k;�]l*h�8���ݐ�}�8�S��E��}>��2�P���ɷ��4mlD �&xI}{l��4��b*{?�́w@x���֫�o�$����4�#*�7)gOP�NL!W��&��g=D g�;&�o�ى��eN8&��7�0�7|LoA@��Z������^O��?�*��!��1Q=h؟z�5��vV���Uȝ�sX��t��o�^2�vL$g��ͯ���D> ��\?�r)Dԭ����O����ej��x����H��=iFe;�x���Hb�*�w=l��b�%Anf0&xV�]�n~*�{f�P7�(N�|#�ݲ���p�������u��9^�DL�↗%�.D�j~8U�~�3p{W�h�Se�_}�ޠ1����R��UxFs{���Z�ڑ�=~�LLi���9ʆ2�k6���S���E�I'��I,%Z���4�&�~f��ɳx{kch/r�Xz��u���ٱ߭�h{R�"��<Û 9��wL-�lʹj�!��ϻ�ej���v6b�n]�\d�j\=�p%��2T��W_���2�<"�r\ڮ�>}v[����7�N�)���)��l��4�6Tʑ�*���D���2e����Q��������~:lg[����ήQ�iu/sD�<+&�8�瀚��A��4��8}NX໑�-6
���+V�lʆ'EO��`k�*�/���-'�2k�pd�hV�@��`��h��7����%�)=7�����aȐ�W�qP�R��H��-�|�B$��i5��af��e��K�s����'�y���* Q��#�$Q��;��^����� n˭Qܓ������y7��	�ZK�'cIgq5CE*����=Ꟁ���O�s�[�8M�x$2j`eE�;���Y^���
�����e�֛m3r-r�+i����C>�ؐ�=�ݽ����?C�b�t�(��Jە�s�M��@�s��8�m�(	H^��,3=��8��c#Uђ^�.��^mꋹF�gQ� ����8P�q+��Y���nP�Z�9>)P�n�PE�+��hU� ���52c�l@��E�W�o뤿ա�R�f·^�<2����m~��]�=�}(^+�/x��!���N@�SS�섗
F�`Cm(di�l��/2�� ���y�q�ʃ�h�ˢt�bg��5˦I��K�Q;m�6Q�B�����E^#�Xf[a��)�c�G]ӌA9���&&ݯ���	vFb��9
$��@��&]<p�-��2.�ԑfp��6l�i�Jp�I*r��I�^WX�7��j���Oj��<�	��/n�1�H�1������ܰh��Q�'���pmO\\Q�'�ލ��5�i�!�js��0>p�0/�A���	�)�m&L��&U��7�����W��?�LK�-q�?��rL.o4�С�W�f�X�|�\�������F�ىC��?\��Qd���ޣ���N��:$.P����L��ZM<�����d��dR��aFm������Z ���/xڙ�y��{VgK����9=sI�jH��|ϲ4�#毦��}0[_ո���'���v@T�*�s&��K��_�Xw,�U$FJDh
��_gjǨ5d�����o�6���j��M�L�VN�х:F����\�0������zm&f� F�Ӟ��0����`��<�Q�,J�5*��F1����bz�:u�@dq5^�`��f�^1;�R
�\�^ ���u����z��@c����z=;++Xy��[�F9o�ٚ5�l��e}ӏc�ȭ:����CJ�0$��>h���`��� Y\�QZ|.|F�=z�Â�L8���d~�A5��w��J�z�HI����B �`��&CKt���!���HfKZ̺�)JR��2URK7���3�X�Y���pG��ʥb�Zg�Vܐl���c���1�G� u�Q��-���Kx'ϟ�^��J��1:D�%��$TIOIim�2���k�#6!S�-�Q�տV�n~��*���`S4��ס��D!���mɡ	�ٻ4%P�W�%]ąh̔CS���Z;:�z���"�������xuJ2^�؜��r�ɗ=!�!/�f�=��nR@l�uL'X�6ȭj�_��w^��d���5����(��`�ø���P���*1*U�����Lq-/��g[P�8cϴ��	7Ƭ`O�E�G��#r7lw�r����+ڙ[��������52��i����lAQ�v�-�%��񊲍�b6k��[�-��!I|�|���5zZ���к���(j����0�M�cbP	�8<_}��k�.Y�<w�B0G�GH���?����z,��0l�S��3%/��E: �(��y&XI��Қ�Z_aG��!K�L�JP�]/�k����������ɳS��F���� ވ�r��t�s��Р�	;^VԊ|�C�m�D#�?\�繹�D����nGED��6/�h�wf����gs$E�J/m�?��_�c��\�[x;�MrIz�Hg��yZ�� �3��L+[��Җ�cT��+}�_,�*��(nn�v��ɨR+n��Xz�l>��������ˋ�9�-���!�>=�&�fY��r��l��s��"^���W^��zp`]��7��*�����H"W�gz�Xg�7�~L-���q�{�?��z*� �v.ռ���d�۬0P{޳�������M�&��l�����a/	G�K�G�wd��cK;C��#��NP���뚍�݂���[G8�s�N'��+G������s̤�m����{B�?�t�?%��K�<�.EzR�.M��|�ŞԂ+��-� �dE�2�m#����4W��J:�II� rv��C+��q�]d�YG0����U���ڲ��,��/8`$��"c��}1._{V�����u��-���|N�\*��To�bd�A����5�I��99ܔŒ��Rh�ˑ�}{�?���g��/md��A�	�B��l���L�Q3�t�M��6��������mtmC+H��Ѐ�'p��ʱMW���Ug�љI���*�k�1�z��O��a�ֵ��S��/"�:�aK៬���,'�}~X\��W�Wm�����zJ��5ק��y�O3X��s�YZ��@��C�:�����oU��4�H{aCڢ,+/�R�G�߱�������\B�H��5�IS�:�g���^��8	Zk�S�O�`֗�z�$�����ٲxe��w���^��rI�;v�g�D�0T��Y�a�D��꾋�uE��"F3?eE�PSOeЩ�6��3�7a&��(�Z5���m�d��u���p����:8��k|6f7.,R�S9|���l bW���9	NOm�M>��Ih�lGn�I�;�稶�o���i��c�3Z ���=��\;I.��S&!��!����'!��Af����窫��fY�Y�`)J���y��/�<�P^p��n����.ZT�?�a�b��UŁ�`;��e��,ˣh�B��S���{}�q+��'ٍq�X������U�kJx�IG�������_�4s������w� BT(�Y7��	j+�B+��}rz��� PdEC9	���ڄ}��XA�	
�Iȝ[N��� c@��a�M��_E]�)[
�[_ j7�8>1G�<�n�.˛���5Y�Fn�!�g,�^y��y�e�p�����;��`|��ޕVW�+	��oOnk��C��K+g�+��@���P��Lv����~�k渑5\$%5�V�*��'i�1�ƛǵW���0t��9�#űcX�����VХ��D j7���d�O����BN��TW���"���$0D(��:��P-^�0dq����г�s�Pͽ������ E��a�P�w�*Ls�з����?�V���F�'9ͥ� <U��߇�7ӯ��q�.<������=�ц�4�  �(�qU�|���;��P\�T�d#1F�z|{���,2�f-��A}�*`K+��cك���_=9� E?!����!��q���,$tlaҹM1ԧ_�hp5FV�[�u�=O���3�������NG�#��������T���饨X��[g$J��V��)��YW>'Μ����|{$�XIPM�դŖ�u�Y�W�'ێHs��y�J�}w��r���>���EPˣB��Lm��mq0me�q��&��4��N���d�)���Y�؉��2��! c%����b*U����	������ؽ��w�t�?����cGᇐNP7N��c����Hә�>�7vO��1�38�滗M煘������iDE�[)��`F�k�w��A��	�{v<�zդ;-$�-��j��#L���uT��RH�)�W޻I]@U�:�&�~�I��r0�q8ڦ`۽e������A�۵�E��8��[����x�$�XY��x�]���s&ԝጁ�e�>���+>��Rm�&�h��}D6�U��?�Pnz�	��c��9����%2s��v��v�)��DI�l!"����#gӨ�����Y���1�%f��[��������	�s(��c�'B�M�_����wX7�;{��	���'�x��#W��N1'Dc?���϶;��0����G��n��L��I�\@e�M%%��M���	�0� �X�mG߼�0�|�t�ޯ����	AH�U��0�n�T�xIT����-7�o����'j���Fp���M����\2�RzIc^�Y�l��9J�@�L����י��ܜ�0���~�|Є `͠梿db�>Dq�t����G�v��(%ؔ�6m����TU�GE� 
�ә4���H��ϣL�u�ee�����Na�(�C���$�M#�������夀#!&>�C�r7Dz/鲎,уl���%�L=O�p�+A���%g�.�3s�Ys/:��-���`1�{6�����u���`�}��;U��9��5m=+,�fS�:���q��hk0 R��7�u�ai!��҉b��("���6H�h�+:��-�dÃ%�O?g��>�&��z�9UڤZZle�q�a~�ـ����:'��t(<Y�nlD�1�JZ*�hL�m���G5�p.łi!���}��_�q�J��8���NO��-�N&�¢�Z�4<wF����N��+,ٱx��/���ddj��u�W�ף��.��ğ�q�+��r�Cw4M�Ը68F�`�#�Fzu��W���vU�i��O�Ɇ�;[E��
�H� D�J�z/�s��.�)�yp�ې\��|�!������'˷�Y�~�o��ޝ��<�����75�p"	sBV���"0��	�vl�N�h٢�@�����П�u��fc ���m�ti��ҕ�9򎌍gVp�<眊�m��2FȖ�A7�
��4��v��ESf�4=F��d�nZ@��¸;�ϤL�E�ȅ��\M<6���fς1�f�Q�3 k�ޯ[�B;�U�'&�1�4_�
e�0�ؤ]nzc����l�&���-R�^�,��T�gcB��*�pe"xW�L U�E���i;�(1��y6�uj@�-%�K,��=Wo9i��5�u	���3U|�~���A�h-Gp��'s����P��d���Qg�KΒ��7�^�Z����؇֌wJ$:_@-����������p�{p~���d�u��hi���ou�<߇�^�c��o�q�r$�@I+���.*�����y�y=Lo�w�k{��?�/9��1�7&#��v��5'氍�:垮n R{�aH�;*�B@f	b���I�ӂ���E�)��J���Ԉܛ��=V��  �Aش�X#M�Z3�9g�����]�42!q�_�A��hM�w>�Q����:��v$�U���M�eM-�_-]��f�\`�fJ�K���<��ųI7� i`�%
�M2䘬ka�V�LF$Z���b�I��.i}�͘�I �K
}�kr�nԈ�I0���]��q���&o���3����!���ن�@��ԃ
E�8��`�)��;���T�����RR�s*
�7��v)Z��3�y�Ah���;
(-���y�=��kD,�`����:zf�e��Y�%�323BR5�}p	l=��޵����P@�2�v���O3|t(	�%9�p�~G�5��q�����_��<Ը>�K�T�k�B�+���c����k\���h)n�8���?V8�n�x5��`~Ƽ`�x �Z@S�b�4mz'J�wh����ڒ�N��ϛ��y�A�����v[�����Ў �z3�pe]�r	��'�	`�Jp������w�/���Bx� ����=�Xn+��%��>_Yv>3e	��� ��n�E�8X&���*�>��$��Ѭ]޲���aK"LsGl'lp���tq3:/�ڔE!�k*CAШ�yY�&�t�62���|��H�iT*�E(/�r@1sƦzt����P���R����:���jO��a Ӓ�b�\ds���V�z�D���eW�T�[�b�3�F�ovP��J #s���v�->��p�ܖV��1N:St�H�Y�z�xBZe��?=n�6hp��#�\��i����V�U
�����`��*8P������V��vGY�� ���2G) /-�y��9�.
�#��������`�k��i�_��Ȧ]L��^_�,�Ӧ��8��c���DB˙q�pޥd ��4�����l��=�Y^���{��s}tɺ�\�;�oDγ��8��`���=�x�A��>����g�p+����2���Hv�5?T1�0y��.)Qv��E���D��eO���0+7��<0�R���"9�h�ơ�1���r҈��|m��F$�l��N�f�GՏ26�I���I�&*JUs<
 iT��_'��E
�vr[��,,t��*�
i{
��_��*��vM���J��ͻSP���<%	��&5�w7�"<�G�9�<M�ݻ�)!�W��16[�&*��N�}����Jq��l�|��Uj	��I����juJbߋ�,WP��i����A���0,�- �)����ASmBh���?���r2��E�z���:UT�pe�W{�DhI8�f��)���HO���I-5"��ڢd�iP(�V��N�ئ�����J��;R�s��m�J��H���@�n;�����PS��>�`(��F����0�������x��6�P��i�����Š�%� ���W��Ϫromi(ŬI%b{z���Q~�*�3�7ū�O�;��u�����ڌ�b��P\���T�V�.�R��4�<����UY/K���d�%��+�H�R�\��Zǯ��X�a{lL-[�L`�����=5"�w����/�R(V�={�)ǖ�c�4n�i�("_�O��px�V������d.����C_|��7�(��U/g}�5�	Ǳ���
�՚5�w*�'�B�'��5��"%v�!��'�*����H�nB�.?�������J(`1/�]8�=ŗ��Z��'(����𖄭���eް�Ϗ>�GNb�"�=��G���P�.X~7�!b�kHG�˭�GV�=�"�Eo�t���7��a�%�Yh�����a�i&���{b;�$���U*������vh���2b��Y��_��+��`yi�a��a�'�p_G,@��t�����&��7��[�H�їi�Z�2��;<.8��7C'ߞ2�@�[���x�b<��#�Q琇�i	��ל��&��>8����9��b�Ë��wNmm��u���\/�[�[
��b�:qZ|�ކӈ;;.t{��k1;-(ˤ��������F[�C�b���UtE.x*��.#��%}57��N�k��f'R�οB;?$��>��δ�ƨeK�1g�ߜˍ�D�u��cl�5ހ�f⇨\2OY� ��K�{��7�i�!w���hlc��Y0�~�h0H�[����9��������%S�� ,��	�$0�y�,<#�ںE`�W�r�vD������4��q�o�$0�����_$�ۡ.}��⿘_��X}3���^�_m�D�kT�Z�m�,[1�ĞW���Q�zohw���VNI��^���$N�+��]>��5�_X�<�@(I���1�����۔ߪ	v�Ie��ΡJx��3��,Ō��������a�p8�����։�5u 	�An���K sR�qK��P����6ܤ�iv?��2�T��hRr`S��9�d�cn���ɢ�d��,  Үm'�9�v��~p� N��vL!ny>�dq�B�&'=1������s�Sx��ˁ���E�H�A`�e"/@V����B�<�����!��	��t�)�ՠ��׸��~���Q��y@��\9v��^���-����.C��mw't~�^�-Ӟx�F�2L��r[#2���� y�^5��s�@�W��ZEm��J����L���$?!��*r���z�y�Ykd&Zeͨ�xgp��b���q�T]�����-�X𔨰�/Eތ`��
�&]�6�D��{B�2��mx��_:��:%����2�_�@�all�j��� k�#B&����~�G���Y�����+�pvirkI�>m%�j�����N�U�bL44�gk�V���z�͎�(_91dZ���|�8QN��*pȣ�n3��N��Y�+�� �'��Lb��?�$
pP�+��o� �J�9��U��os9Z�#Ï��l|SK�ά�:a�۞��!�|{"��������p�S�����$����@��A����V��t�1�c����;]�'պ�X�t<Y���چȲ�~F��UODz9h�H�ᩖ�J<�[dt���}-'=�$�1� @�X�FIv��P&J�	������%�rU���07%L0��ϟ���S��(����r� ���J`�:T����';�9��Rp�_ b� Ȳ�{/��6���z���V��
� �k�%*�K ��<F���`�qs���v���!�K�����ȁop�B���,�����d��ޭX�f��b��H]��������o�:����
��q��q����ū�!r�^V��<�?X»w<���I��<�`O�Q�!���ZG��r�����'��Ľ"�W@D
休HeŃ�T7z^Eᗭm\qW���]��^��m��<��(���sW�)\�",M�bR6�QN�69��s_z���� 	V{�)i��e���S���o��RC �#vk�z$
��l7E�s`�/�ۻA�&��-�L('*�$pPD=���s�:%<l��W]U�Joz�ϝ�U�&��4�"X���.Bs�U�����+0�jygߺ16<(�Z�n�T����>�=['?�B�N���@�s���{��zMP'�ͣ@���M�-��-u7d�W��c��m�E}e۔�m�q�D.	B�L�Xxa�I�XE�G�ɟ�kOPuE�`�y.#�����A���eKMC���+���e�&��tޥJ W�g�zF�����Ȇ s�2K~��V�ꇼw��Sࡓ�Ǿi�Ŭ{�}��S�R���{g�+�*�4J��W�K�x�ߔyf�U���r'LG�
ꮡtҊ�2��@�N�i�_9l�;��Igk�����z�|eD���%l��ծN�n�!��+�v�	����E��C3R��c�{�
!��}��B�0FӉ�T��n?�ō1��L���o3��	��G��x������5���Bw�l.ĸ�<MZ'7S��<p���Lt�:H(d��X$�'p�v��7�� �p�#Т��a���ƌ�J���S�X&nk1 -EkO�HSM8G����\����i�DP=��I��p$����d=���9u���	]��w���]@�vC�hK��:wx+�" �Ι�������"$d&�
\I5d���~�� MG�̥YW��p�[V���59�X�=&Eqx彀S�˃Qk¥��S 2�b�����qu�f�@��<GSc������}�,ݼ���x���Mา?��E�|��t���q�@Z>���~r$ۆ�d�X�G	�d
^��hD��z��cM�T_Q}��l1[F/-z|�G?�m6��_�Z��F�p�B8��,�Qp�e��,PJ�襭���MU?�����[�!O�Y e^a���$щ�^v�7O�Fu�q�W�w9�#�N1+>�7T�x���)�due���.��c���
�����9s��4=�6��Pu��n�hrN���ս~H%n��{���&�=v)4���v�T`Y3�>$ݏBxs����K^ɪ!����z�����W缠�l�e�vJ�&�ld�(�U�U�y�(���Mƺ������$���4�){E���Q$�4#M���`����
q5�9���\�f��8(��l������AX�c�*��R��Xk��%����u�Uu�p5��͖�n{��ǌ���_��v���?3�k�񁬆� ���t��г�QN��o�۹����6u
-c�����Ww�s����h}��J�WFʜ�~ѝ�aU�jp[�c�֯��'��B�,���9�X��c23��k�|�Lv8���-sx}��������h�ٹ3�Uw	"���k�B.�75Mׄ?�a��T�8��]�k@�����CI�R���o�E-��w��zt%!��������o�C�&�Ti��6vx�7Q���K�\"���v��9�t�u^e�(+�z���ArH��9����?���y�&|��4=m*����C|�	J���|�qX4��216��f��0�q�˷�����H�������L�i�Bl>�~�+ē����o�K���g��)K���b��0��$L�w��f���GOޞ֊vH��<R'�T��W�UN�"5ܻ��w����\�9q���!j҂����A�FT��$O%Yg����?o�`��,�&"�J�[�K�zc��D�3\}(%Y����J�2,�Θo(&X���ڣ�R���釃h?f�K4�x~ˈVP��Q�.�w���s[�+��=���am�Ѧ�kLl��&��9O������W.\�Ԁf����XN��8f%�?΢D�ZZ�X1�.hV��8�"YU�ڃ��������@�v��%��Z@j����7,Z�ܡ��z4w��И:��2pu>��
����"/�r
�o ���Z��4���q�?�ix���ͦ45��W��?� R+�3��E��9�Dέ�S,s��R���lD�EM��Y{�6�ZrfHIgd��Z�`'��Sh���Z�N�m�%:N;m!�]%�%I)����~"g���՚N�z��g�F>���W���:���xZׇ0�����*�SZ��M��� ��QL�e�T��lk�v2��$����3Ai�"`ɤ~��Z�Y�I�?��٩�D{���!�7"H-�;�[�$�~+[=-g
�5~�P��^���߱��
{�ji��^y/b�e�+|	�R㗼ɢX^/�v䶏�]�px$
�B%��4#�o�#Ļ�2�h��Y,���R�_P�:�9���"��=er�9B�rJ��_�
�/������5�:WA�t%R�<	�TD]A��oq?n⬴"s����~7�ϧ��*�5���'1X=Z��f�`�"�� �1O0�F<�Uێ�j�#���!p�{���,�r������,3����Mj僇cǰ_5�@3����p��7~��U3����I8����wg�{8�0�y(٠97�^}锹q�a�%/GU��oɠ[MQ���9���sH��Ny&���|e�Ud�����^u�d����G��.����;�_��%�%�(�j4(M��{i{�{�$�������*Kd!8"V�q���a�>O^n��/�dK,x�y��Q�@��y� �0��K���]�Z����@eW���&��˛� ����QA�� �]R|�*���]ZH��qq��8n�v��?*�
�>gN�@ҋ	��xm	:�܉
�3P`���2�����g�+��#�,��P�X�I��":F����#��R�q�%�V>t���ӟ��TcC�Qc��L1����ߚ	�L
��e$��ĊURt�Q����Q���bF63Usk����K?PA��l̫� H��d���}�&�
8W�Tf8P��{�n^(N��Hv�q/�߇��*��S��@�(����.7<�@�s��:�J�Ej9�V�'�Mc	y9�	�|4�O��lH��1�'Y��O\Gѹ�pg����T\���	lR������&����N�f��"�=���ƈU�Yu�n�7[CuxX~`t��FK��RD���Z
�+��)�c���(Ok�v�ܯ����'��d��aRf�'K�P�t�[*�ܩ��� �e������Q(8C T��������u_����pDԷ&�1˶a7��c�"n?�.\�5��A��%l�|�2�@�$�q���jY��Bk`ܕBSs�Nb���N�_FO�=�Z����Dd�l�~�_7��SZѤ��WW>
<Jt��X�I�;���� S#�<\R���ܜuތ���X�S3��zN+o	w��K1%�8�m��ʡ�R�?�� �֢f ���I� �J%�2,A��h(�'�¡/����^�뇍:0se`v�2)���|��!�6?�'~�ҧ�h���B�4�B�� �-���&��xp����$�7�&��wڕ�e,��b<�~+���4�8?o��w���0���B�|(��|�7�P�iɱͤ�̀6E�a�<�w�h]ם��as�^�w�<������U
7��;��HKR�=�|e��h�
:���4��W�qNKu��7v��ʵ��n	������mWri|�0����}{/��b�B�v�).�  E���f.��D
��9�+o@C�j��z7���(��V9*�y78n3YRO�a"����4��_��12��
C��p���j|��{	���A9�����~*7b�g xo���K���O�K�:����l�+�:[~�.�0�kI	n��$˿��'�~��$�Skڬ�)}�������[��a=�N�����u�$�� x�l���@��*1�!b��vv@���j��Uc�����9U6�y7B����Gqg�a�b)A���V?�`^�Y�EǾ_Y�>ʍ��X�cUU��魧��A�p�l@�0��}zoeN��W��H�/KO^��Ͱ�7��"�s5^'�R}�Ƶɤaz�����ў=�RO���e���ye@������8,��<
�?�҈%PAP(��*&-_?��W�97s���V.� �M<��ܧ�$2ZA�����ܗ�U[AI\7F�t��}���lQ��(ώ�n��4o@ $���I~W�^�z�ނ7c샍��ڶ�bB�U��)ԗzz�9JEMY�/2��E�X�B���?��\z����$ރKg}�c)����)��3AN�� �R�o�����轌g��'�������Z[���l�ꗧ;��S�гr�A�ۯ�fe���ҋ� ������E���	R�����D��IҁWh����ho�ϙ�s��=�S�UD2���Q8m�� ���� �HVl��S(�AȂuǿ�]���X|���&�~iW_`��ҙmA�큺� vI^������ĉ�F[�bS���m��C`Ƿ-����_��M�A1������P����DvM�k�YJ��A�����ѷ�+#��۹�o��?
���fĮ�}�Ǐ�������	G
�����n.d���2eS�o�FS�c�^&���E�׼+�6�3]��!l :@ֈ���&�ä���^�`����|�4���ŔۖX�Y����9iP��N5�2Y6�n?�V�0��|�'q��K�b�Q#6�b�:3a���u���@�+�����nCc�t�m�,O���mt�X�9a����+�����i�C9?��
��9j)J���i2ʰ0�Ri�ޮd��E�xs�R5��8P��cV[�M�ݧ�x!6�
�����$�y�lU@��xK$%�S���O[C�T�߆\�B��\��Yx����]�ۇu��W���%R��93���!,�?�О�4c0��4��A�$���3��6iTI�'\���wX���d��V���9���n�5RƯP��g�\:�]_�R7�����t�6wT�i-�]I��=;?���
T�R8w`��_�����1���dEx��ISJ��eI���}��f �,*�G�0�9����q��}�a;�&��?I�b�3�b�ź��0p����҅�V
�]��zz�J�3o����.�\��0�v�2#��w��N�
��C��/3�|Ѐ΍6�j���n�E`�#	�����C�AUdOQ���.��U(�t_�E�E�-�W�Z��el޾:���.s�9��=����>���C���C�-�B(�2��cdZ�� ���+�ٹQ:L�������	�AdŸ�~o$pp���tɻ�Jr�-P�@^�y�6m�N�s\�p,2�UG3K��@��9��~��co������*EX���2uY��T@P���-�EX��f��s*H'�Lv�xx�������:����'�6A|Z	z�fh��W���P��:9�	��5�lmK\}�lX�����v�~�Ky:)Xo�R�_*�\ns���o����v~�1�^h}J�7��$�Xq8�U�i���w�uʥ��3���N�
�n�/hf������WJ�O���u�O�f�e�֝��GVz��'D@�S{�+MT����K��{��A�>�Z���� �1'>�m �2�S��PͮB�/Y󦐹ն������ە`��?V�}�v�'noK:��b����{�V�)�2�)����'�Y?Bm��3��(Эc/&/�﵃-V��^pU;dm٨k>�m\�qSNW�
�i�-�1����ů�b��O����	�h� K_����f��������0#2h�hC9�B�e�yu�V:�g���8�/
mC�>��t�4�\��1�����:�"�d�3��T|e��s�Dk�g��5�t[^��J��KImxr����J���j΋�-f$��4�V|��N���ϋ"�j�v��#"Y���ZE~¡��|=d��(�񡪊�^��ѫ����~�	ϘGU?|����a*r���kK��C����KN��<���v�4��q�J|��\�����Kk�	�&�o�U0R�߮	A�~������i���{z�y^�
g:��IG�]��/Y�&��.���)g�|��o�pb6�_j_�I���Y�y���(�{N%�&�o�)Qjuu��r�'Ϲ1��y�<�:B�m��[b+�*	�4��B�?���l��!fc:1uP=b�Y�-�3��u�U��b�x��X��$!.�4�т�Z�^���}9Z�Ă*�wl2h�^�$�k�{t�"2 ,	�?�~+����Kh��R��wR"ݯ]D��@�_�!w{�o�ީ��,�u3�7��x%�.i���lW�	���4�| ���X�����l~ɔ���4г���2�Bg$1�-�
�b�A���7��ߖ���;&�)M��4M�c�Y'a��ly$�����	Y"N��	Y�۱���u4�
�r�c�U�OÝ���]���ڨBf�i�<f���h0��!�O����N��R'-��I���(�6���re������?��)ތ��N�Ԕ�UB�Qvff�Ɂ����xlW���SU�G��狁H�1ǽ�9���@����~�����"(������d��¶����c���?W���<l�c<���%��r]�Sof �V��E�����3hr�P4�0S�sH�{'� �|t�L�;��:�y8��ӂ�gUH�kD��Z�-2�GlTnt����%2՟��5^�f^<c5��	�.���Ӳ��%)x�~���wp����ٶΧH9���戸����b`diɳ ����2���ȟ7���";��,[38����k݊t�La�J�`y�&o�����|x��?3]a�w��juI�-�$W�Ƅ*�K��[��5�%�3�m{�1�pyI_�A�m�ª/վ��c��${�8�#�3�����aKLjQ��n���_m�l�|6W+;׵��L��x�8?���Δ�쬃�|F�e-}�������6鵻�	wj� ��E�v��۴+��p�|��H��o҇e�JDz�r��OkG��MA�Ի��/�9������~��q�r<��o��:�ӅҊv�b9q�����khŠ�ӼXl���uK�"��f6)��L�z�@��-o�Dj�趉��Nx6�zrW�.����}>+����V�56��mwv��D��0��[�O,�_�A��Ӹ2�f�UQ�nH�]|�IA�m�X<�~%v��@�7b��$x�O=)����\T)����i� <��B���(�:j�Y�Z
�8$%;�::�׺���_xCҟ�v.)�j6󚻽�T��\xԃ�8���Y����=@����fyN\Ş<�O�t_MW4y4"-��-�`n~�T ��<:*���k>���<fC�|:!J1U����/�{��S[����I>�q�O�+-��z+��Aw�#��8��S�1o�`ѱ�%�HČ�q<;�tx�c��so����|"\�����QCL?`Em\� �&��H�1�o�%�=�#�uxKR,6C~�"ul���������Pʠ����LkCCn��k��6��z��dm�P�d��X��X���״�G��3u�������6�4�P��mEܶ����\���ĳ���x�1�M�N������.�A�2��
���nk�+�� ��i�,���?o�}�[3)��+�&��ȱ�8nm�N��d��M�R-�Z.�̡��F���[��������H��ޖ7!Ȫ��`7%\����������o�5�����I_B�s�{�FB�3� ��i�B'����$�Yj\?Ϯ�C�����2(�gAj��>���������ݱ�shʁbLd\=�0GvEr4	��z�fK��U�d���Iެ����K%���u�ژ'6Y,z	��Gkq�&��&��ҭ�����?����U��OU�Bo���g��nhxh�^���	eTVh>�<��f��TZQ�$o�{�h���|���do{�N������z���O�<��(gg}+���M�D�d*��69�o[�!k��7�gBfq��y����M�|~Y�
W���� -��]$@j$PLe��@�F�aW�e����K���?�,ZL�.�(��C�/�fH31�7<�33&#������Ku�@�ƹ*��B#T����Ox��ItdY��b��]G�*Q{î�&�}ϟ��EQ���TV��~�׀�B;f��#��.�y���O�����2ۊy����B��V�ɪ�k\|�	a��P���l{Z�R��dl;V�PTY����1�� P�����CC��=�^g��ϋ�jj��LQh���53�):�1����9�>'mH챓���͓��#N�)��\�&2����Հ�]6�3�O�ı��
��o�4���ߚ稛��*;ߚ����t�P��.��8��Qi�Ta�+0p����/E4��b���y#;5 [j��(��*�I�u�!�ٝU� ^�<�i$q�����ڡ5���${��rkՑ�7l�a��MD}	�'gJL90���v�V��/�|@O
,4:QPynL̑f��#��v^'g��;�l�Ӕ&{-��\L�T�
B}6+��Ȩb'	���Ӗێ0���p<dw+��N���t����܈�H�M̞���WS����1^�?�{�@�i;���P/__O>������\�p�S��<t�Z��L�-s�+W��@*WS��S�374��Qk,Tڈ��
�a��bD�� /fi�EN�����GH_c��������er7!`VF���������g+C"��u}#�X�H���E��_�"����S���+�	{�>��Ņ��,���a�g�̒\��Exl��g�g�s��6��A��يڄ�}(R��I���%L�˰]��W��შ�E��ф 3S�f�,t�xu��� ���K`���!�Ξ.`
�CoP�b�Q���>^�G`��q�8NR��ǰ5q�H��#����{��Ӫ;��@�Ói-�B
�6��,SQ=�7yx⋙#�Ŭ�R��FF���]��æ)dO�G7��t]�$K'�r/����U�O�E�+�'��������wdi��9As��^#��u���eGڽ�`���ʮH<�а2��M4`f+C ��a� "���kǙ�����~K��U�x�fp�����7�l���a�V��yF�f�)���G��4���ݚ���c	:��*A�'�|R��*�r<�����o@���--c^}%d� 3Zd�Fz���S�ѡ����?�ʻܷ��fYw�k¡�q�i����M�4�Z.ŀ\]W�s���Oۂv����u`s�a���U�nC6L�?� ���P�3��0��kVl��z#Ap�j�d�D|�<� ���[�#�S(��>�g���5!��g�(5�k���z�,�c�������ו�S��UJ�ӗ<�Г�oze�]VO��q���_I��.b��c��뢰�*>.�$q\>Y�n�
\�������(�P��~B0��#�a��K�9N��*L�U���y(Xm� �7�J��@ՙl��n�cJ�U��ڮ?�s9���ѽ�<�ԥ����AYwB(��:�����H�+�U�=�e�d������z�dX�������!{�pMA"�^� �ca��� 3ۚŨ�aO�I����|��zdUc�s�G^+kM-�V|xy��SN&7fCd�Tq�۱tP,��Jb]k�џKX�Wo$ 3���%��i9M�K��Y���ߤY�����d�nI�e<M{l��Q���S����т~�I+�pm��`%(G+@#�t�7E+�H�,�%C�h��U��]φ��_��_����'����%�r8�1qp��S��ȋd�{C쒥>���t�^|��V(�_�9T�a9G��`�*:wg?�90k�u·�63)��E%�ʀ>����pd�E�"�K�c�7�*�9$�S��,��Pj�W0@�%�!~�~�G&W	�{����d�1pJH#[��x��IRF������vI�q
4hp
~�9���.CW���#��}�G�	�a�����L/�_XʹTmx��M� \�p�"���E�3/]��%:9b�v�u�k!���,ZkN�D1�Y���eչ�R(�������ۣ�|9\�x޴�$�=�b��SDH��3�<�1��E����~WK�����:e�b����s��k�aZ_��P?ixT�G�l�����X��#u�����:|ĕ[u�:��� 4Ռ�Hn ן3\�����̮	�9�Ɇ
�=>޾+���&��r���D�����%�8��:�3�jCv���8�|ȵk�휮P8Pώl�[z��Q���pŲ��Lo�Ky���>MCu:  v�T=�N%���a#Q
��
�I���L_/�&����fM`���V�j��`���/`�!����_�O��{6C�&1T�Ơ;ɺ1Gн
W�tt��>���
K�I[m���J���=�w��u�Ѿz/�-�P�˔�'��~�|���������_��$�Ϫ�*�5��� �}����{�?Do�I�O�̽E�2kB�Xr���F�ްT�����s��P�PF�6A�<.O���
��ۏ�dSy�%�,��k�X�R���[��y>͙�����n(��A�_K�1Iђ��r/9u��'�g\��e���|Uq�\�iuA�*�vCVbW�x���"s������$/�&!Z�V���96%I�i�'�ex�35N� ��c@��K_t�w>`R�e�|؊Z�/=�mT׾�"O��vs��B�m���B2�>�!��z���zJ�T��wf�ҕM�d��Z��5*���t�-P������ ��g*����i_E0:�H���2�i&<��N
�F�1y��![*���7���a<)�Jm�`T�
��%~D��o+r�Bb�M�>B� 6>K?��3*ӭ �L��?cs>��%D�g��t��>+� �u2`��{�\�x�"�o��2*��/o]��;��Z���WR�e���"ɗ�-�9�M�؄��"(9���ˋIc���c0ܰ��	1BC�0�W
iA�'�k�
gO-�=s=��`�N�����\pkG�L��I"{��?0����/��/���	ѓ�#c_e�����_��s(i/�$-ܒ��;�r`�~�v��f�>�^Y�BB�s^��q�����";]v>FD=e*��4��i|�G��@VXZx�_������a;)��b?/h���?�UF�Q�\� -'�F �;S��!�e�ʪ�w��%��&��	h��"��g��%��~g���<,ћ�LXC4
���������(H� �C�}�>��k\���;��9h���Нka�y�A��"��*�!k�ªv �.V�k��t��ڸ���ZhJֱbd�]-�fQ��[���WMVg�)��o�&R�X��c<S�i1�^���Q�M��6��d�Q�Q�-+��}L�{a��t�L2���?�r)���Pށ�6i/V�.�'�Ea:1طq�c�#��+�ʠ�Q�]`��5�S
Gu�Q��.�/�8��j��W�z���ir̷U��#+9bKn������eٕo"k*�w�+N�xqh���=��ǬV��?wd�Ĵ�����^3\a���?����'��G98��b
��v��D�[��٫�[
d��m����+�m�P�`��'�ȟd��߁>���UrP �y�WZ-p�w0��L���ӧ�/]7�2�@ɝ_�nA��R7�S��� ��6`�[K9���H���=hGH�����I�ičD�P����ߑ�ߝ[dD��P�,�ȼ*��x>�G+��s"'������Z�ֹ����^��>�h�~T@��*Ql�Lp>���#�@�Z�_�2L�j�i��1>#��J�l�0�Bm9��K�~�gӶI�(.6��5~�G
-�"�#�����D���h��i���7����sLK~���@������dW��)�#��'m���!B��B7���5���l��GLm��]^cZ���N� �xum�L��d���d,��Z%�qXX�%#�	�ڤ����w��L�S�r�j�}����g����-��n��k�g !L��_��^�r%��'�Ĉ��dH���c���]��P����U���ݜ
{*��{n�r�)M鿅�)Z
�osÔ����{�
����.�W^�Rqћ����b�eV*\*Dh3$��V��!��)	�wě���]Yn�\�-�2vo�����C���A������(P���}KZ�%;�D����d�*7��ލ�C�����RU4SS1�\�����1fy!����4�awʽ��o�k��)R�h�|�����,w;��3\�l�t1�4��4�[C-g@���l��G��t�r�_v"��!���&[����{�ă���G,������KWc$���7����IJ
�ǨHI�y�A�3|#�(L�H�Tv�ޮ>�RK����<����ء$��fG��%�냿�Hc��bFy	�?۪6d=M5~D]'��Z7�H8P�ۂ���.��oV3�?x`���) ��ls�/��.�x��O�I���}�A���>�!c�B&�92�`�����)�m���(�=VA �׻�ָ 㖳����NT	HX~�JG}�r�gE�1���k�����QDHM�4��ى۽i�����:�9�l-��á�ۊ��D���'̝��?}��'��'���a��p�x`���+8O��wYNu�;��΄vp��fD[O����E�S��4�Ě�`�u�1(�I���e�-�hU�%O9�u���Aŝ=\bf�+��1US�tm��%"'�|�c�.���UĠMl��3X�u��!��+�t���ظ��QCAbj��:唂�+rM�����2�7�_����]�
bQ���qWY͖����͠���/QϹ[,�N2L}z�{���ܤlT:&/�t�8�7�͖{��Q#}�����;|�Ė7�i�{E�"n�'�$Vk�'cn����K��±��`�~���U�>�T�a��+_�"i\�����n�"y��K��\��;·!��Dd�,v��q�};r�Ґư]������+�m�'�e�$ :D���v�5�јq~�����/�m�r�Tu�ɿgh�i(b�A#p��(��F_�
x-�f�h8���,V�6,l��
���������zz�++4����.�t<7�TS��9���:���m��K��6y���vH(�uW���N(�s���ZQYm6A�<WO=�6ʽ��ѮoO�į�r;��P�]ɱj�Ž�?���!�!M�o��!�;�ݯ������UC���AN������Ν��p�!!,eo���j��M�!�� ���G��xh��O��5Q�sz����?��. &$y�[`?s���js������z��Vߋ��Mu)�8\z����.�䠹���ߋN���=��z��ջ�~�	y#��P�1�<��$
=ގ���S�>E6 =��ʁ=��r�٤�ih�^H��3MB�䋀-)@׈�E��
�p��]V�����ɡ���J�}�}�?x��i|����xN�8��O7���c�M�S����Q�Jy��蝉�o
�����=@��eb����6i�@�(s�K=��9��P���2z��d��S�����{���t������O�^>����V��a�	w�]@��ý�2��G�$�X���UZ[Qշr����(�B^,b)�	Y�-�й��}�tK���A�]���y����J7�=����nM�D�Cm�geSt����!��@Z�V,+�͟��ۇi���� [P��;�a0؅�'��o�I۫	݂.�Ҳ�>rS�Z�:���RU�ޢdD� ��YR��� ���ՁKg�m7�ܵ�<򇿖�[s��/�א8o
@T���51��������
�\�@��j"����2�NA,:���;w�·�~��}ʭ�l7��i~��RL��BE���i�W�HI8N�U"�������<v]�1�� !�"n9ϼ8��⻚�YB��y�a��?\4��⍤�Z�ZB��1E�����w�I�t)��ͼ�m���:�������/�Qdx޼��0�w L+��pd��ؾ�]z9��t"�8{��}��b��5Ԯb"2�쨶�M������it[Z؆*;�2�������.%m*���W��9�j��%ʹ�%��:G1�wB�7�	Tg���(�)�=�?��I����U?�,�\/f�����=hg8���m���� ;�N`O�`�:,�N$��HŢ:˹��I�b�?�M]�G㿍�)�`CI��e-JC7��T��L�5Iٱ�Lncw����3����xy{#W��nL��ўN���4�_ꟗ�Ƹ	i����+�^c����@�����������g 7��Rg��t��zj�A�/#i�1U��7�,ƻo��k�a�b��+�Q��y	��������]o�a����g�iS�.玡&����ߺ�:h���F�u���?q�-�8�S&Z�t.jU���qM�����'WfG?"��m��&��MQ?�9�ķZ�I�~���8(���Y�ɕ�(�#}�2=��艤�&n��x��	{dm�,WR��B؄
N�4Ng4Ԉ>�t�$��<�zR�+��M= l��W�(��۫Eq8�|������Z��
e6���y0|Cfrj/ᬐ�j ��L����SIc"����V��<�ڀ�[������Ofʔ���|��+�"�כl���X".?�L[K��$ZK/�/�啁?z�?�MV�a� q8x�z_�B���b_��>*�m~�.��L��6���,�~��s��<���	1����Yr�� q\���\ŭ� ����&\��:����<��^{�$��*�y�2�u��c����Ge�:s����I��#�B&����m�Q���W���(�ª�I�ge�ι{^�����TC��%g8$7��3.��<Ц#n];�?&��T�.�� ݤ�	W�F��ڢ��_�ub����%������I7&c��&�R2�*�]|�������Ie�.VI�l���p#�������hB����ޡ�!�э�[�?�cu�<�]Y�6���EX�s�m�1��'���QZ&qi���6B�_|^A�M��:��xѭePUv�a��:���9DpGr��4`_��,�̼�hko'��u~Gx�
eHb�==s��h���$r_�oF:X���Ά��`�h���3����u��!��P�$�Lwz����T	7�#��,SHY�ڴ\kD�W�ۤ����N9X�O��^��k��������1JDBq���c��v�̾@���'}\x��b�װq���t{�+96�2p������{�x���N�f%.��������1 T��S��h"���m���!��12!1@�N�"��խ�W���|I� r���B%4Ȩ�Q���!�˷�4�S��,�*�{�r���&E�5  ��ߍ
�I*�#���X5�e-��` �R䋢���}��h�����-ߢ�O�g"�Eq�Q�%˵�Y�xWj�zHזe�+;?��up��&��+n��żǚRW�hF2�μ�pǃ�#wۚ�RW훟��-����<�Z9<|ṩ-��}wl�(�#0�b�y����Dz��GD), �^�e%hP�|\ 8���?��aw�~/���SP�{��2�渕2%RӄR��"�4���<]���)���=���v��1��Iu.�Ϥ�v�����ѣZ�����Y���B �I�����w>$w�;����k�-+�������zߡ̓}�X������H�Ǽ�(��V���2ҏC�
F����y��64Iӑg��8&���S���8^j}`7H�K��6�@�_KHŕ��?�C�]y���	'�Hѐ�.����?�
^�,i�H�֌��zR2�O�N������X�Z������W��c���|�K�I�YM�@�)S̸�_v��ٲ��K��x:�����i�;Ԃ���ҫ]w �įH��t��&� ��V�Ѐ���#����uL���&�S"����+�{��m�#�Օ�Ŋ�d�=.5*�5�$s�Ӊ�:M)2`���T������}��/FC�oV{��*3�Q;Ñ<�f^�w�+�i�Ӂ�w�&�9��x����6+)��2�����.�{B��9OngUx�g��a�Ĝ���@`���H��,�,9?p��P*�o����22�6F��z�*4�ݑ��w�o"���y�ݫq�Xd{K���47"��{,]���8m#\)3>AVHo�U�j�1��2Ʃy�{��g{˺t�ƪX�b������r�!=�PX���	Aߠ�f�z�09�sn�lc���?��'�vn�gf�u~�7�"��_G�$��ro<Y��ڽ�r� !�>jA�F����05`�4�T,�aA�deC�N��Õ�Ҝ�� =�b�b��t���ڞ}�wzĊ�����:���"n�7N���z0͊���U(zn�z�)ԘZ���aBU��sX�' ���fi�t����v? :��U!����6aT��5�q2��̒+��W�QsIP.n�aUm�k�D&`C;E!>�s�9:�h1���=��e�|!�y��w���f���5\�`�#E�
P�͖�q��ʯ�Ґ*�?�۫��7�'��ׁ]_ܯ�q�zL	���Clpi˒ܫ��1P�\��-�B����ŷZ���5=��"�`(��shG6���������\��N�I7p"�H����z/�]F[�΢�/�z�eԈ"�,ѕRRQ��} v�Dn�<�5����B}�T��Vs���Y��/�^[�nܞu]�*�!�8\^�(�pԿ�Zhl�?-Q�Hp��|xDD������
�I/�,|�{�O�>I��o��tD���7����QM?${�+D4�c_������}UW�$}�Kvۤ�V�v,�(�!��w�^%}�t�hѭk�jeRw��9�h��^�\xi
^�L�3%�dpxP��|�+�+	 ��b��4"��m0�j�8r�O쐞1n�K[�rZ�&e+�`����Q-p�����m����#���T|�HY�1��3������ྚމ�ǄwO�Hp�?Q�N�faӒiiwyR�s�����%�7���7㉛7C���< [�,~w���QL�-V��!zx�a�^�0�`.u�c��C����^�q���G����E�� d�+��l�*&����#���|'�р%.3ߝ�UIT�)���u�=@.���~(ҹ
��׭H����j� �r��\���������� ��J��t%��3�sʗL��S~r�zÐ	�¦۞$�p>y3�a�_��k��Uf���=F�M�3�!�J"��ɞ$���٫�h�������Xɡq�,�[?s5�G��/��:�͂6=}0˂ʫ�1}��e�%}@C}��p=�6l���$�b����Wy� ���h�!����'x����NG��'���j�dXk6iA &��=�ug��L�N�b}9��?'�V�I��0n�����K����4��B�)ѩ�L7}���m��~�sRޯ���bTC0�o���+��#��35h>���	�χ��E�e�{������s2�\��I���^:��#���h�يr��X�Nx�+L�0�܁��3����s����r���ChﴴI���&��=-�
�t��Z��L��u6��&�7����%=4B���2i�F��D��T�ǥ#�
u��˟�hSM�k��=gs�����~��=MI �N���R5<�1�L��?if��Q��Gʇ@]��P�Gag��ƻ����d���4�EcuV' � �y:��"���/b�-���
�)^R�[C�q����$+GOhQA��#&��Q��{T��=��xN���@��H1�%����qHkf<��T]�mr�ꗶ�uCDnx�?
������7����А�})�<sը��{������e�Ӹο��,r���YޙT3�w?)����b�ߘ��E��K�c=���>`_��!=mq��7AX�_�<��-��ݑ�V��zh8$���~�x�����7؝��τXy;>��p�R��TUފ�P����S#��M|���Η�`��'J�j-��%$�x�!�M�׿n����.�93�xPM��P�H�!��՞� /'k4��|:��6���a��T.��eP8>��"8�;�<.�*3��9��sg��ـ�� [�/լ����M��9�k�� L������/����ز���ԁ��Z%(�x��}�6AA���1r�����u��b�<w^����^�g��c��H^Pz@��M8D�x�| HñE�� <�WwV��5f��C�+����a4���(X��*]�޸�4��|[�I�c
�6Dw薧P)G~_b��K\Aa���`�%����+m쎌�-]:�Y
Ƕ�D�s�m�P�sQ�ũ�:](N�'�]��|�[�r�c�\є��+�M���ݴ͒@�c�4ԻT�T��0f�pd�8�[z���roc(qr7��<��!��K����prRZ�V�,*V|��S0줂?g�I+�
��w�{&��r�^B+J��t\�����c0d�uyz��)��ӧ��;[vR���8��Đ�2�� R�2��b5�(PP6��I�N��j��ً�����Q��U�m�x���ts�*m�N��?ҸVF1�0,;|�v!��<��q��N�Fh`{���ì^���
�0���0�����z@�9С��z�z��A�]ZɆ@B��	_)^��c�)i�@�um�S�C�_o��~����Ҷ���reO�@�gՕ��פ"�e�x<����Q�k�Y�t��
zF PT
h�9�ï��?2V���~�����-1@M�#	�y6��>��f�R� s�^�9M|�e?�!ѓd��w ��>V��)i
)����}��Ʒ\de誱�B��V�����m�]��=S遞�ˆ��W}t���C?�B��>ڃ�,!a�+��(R}�X����qލ��o�� Q-VrD�nƧϴ�|�]������o������Y2�2�0�������e2�֠kX{����t ���݊xd�g��~7α��V��@Mg
s(�&K�����g/����[�m��y0W���3���E�ε�4�L9l/� 3�^?3`��Etb(ۮ������`c ���_�huY+?g?uK�M�#��3_��� �^ң2U�<d�"�����7'������=�Z���K[Q�O�z?\����~����5���\���/�/q���И^# O��_X���	U�#�!�tKwNr�wT�vzOt6U�r
{�s�a$�u�WR�r�|N4[��|�o��ߍ�Ժ�r����t^X4�ۈ���⾟;f�A�_1}�M�]��F�i�oOWF���h����?&�����$z�S>+�I���OŰ���Jf�]�0Q�:�p�1�=�s1��l�0�Bj�#�>�R�2��=��G��b���"άm߅�����q���P�58i�u�/��=FD1#��x'<�1�&�F-�]�;#�&�����E�&v�
֨$��j=9)|k6w��K�`�n�2t{炙�f1�jc�M,�Jڜ�U����vv��ǚ��ٲ{<��В���Ը�^ovr�����	 �ً8!����v̗*�|�[�\������Z�Q�S�u�̅�f��a.`���v�� 2d2,�pk;� �6ץ�p٣���7��`��Mٻ�du�/J�
fQ��6GJ!��<�CO0<��k6;1�7�d�_�GX�#�7�n�F��tW�$���M0�'���5r�--��DX��riU+����g�F��IBڀ�F/�:+��T�EY��܋��g�jq����?�F���2,�:�<��U�q���uv}����}�!��ang�Q8�X5[�]��E��j��˫�ш�%�\�=i���L�v&�W5|N�1�-��&r��YzN�\_~��K��/�W�K��X�
cL��;�v��W%�s��&��� Hwc>��GV8w��0�g����1��9��|��`z��-�_B-[���"�.��f�a��Q�K��ќN����g���qܱ&�#��yPׂE���*�NQ'�j� E`U�j��d�O�p��Lp"�ش��CY�w��x�&C+g�-Qd�t$��X;�g� ��J/����^w�/�Rm
\�=�{��?��}�z�����1ށ�_*��M|�����,��)s���O��o�gj�P��:�憉¥:���NZ�����X�,�J�B��G!!�ƴ"\� ��hE���)�u����H��#~eS�PX��e��t�H�Fct���6��|��dP�|;��LP�:��=�H��9Y5T�Ş���K����y��xYy�qG����Ϗ����e�Pg��'�n��i�b@1�A�;��H)mR�]�.��A�b��(�}�FrKT���ƽBGtnܕ! ��6���CÌ��rPo`j<�]���o��aW����� �W�~޵�'7�5B����`c�9�楣��JS��E�:��<����Tmy�<�6]��raD�wU�3�qk�Zfρ��?z�A����O�v��]|�!�{|	۠C8Z6�筱����c��b/w�hR�N`�?�����ڊ>wh�zTV)kʮ�.]�S{���M��e�� c�q܌��"}#�uyRg�D0C	w�b���To�ؙ���)Uj ��v�s[��|pG7�Xc*s�(Zy�`U_3@��:N������I�_>j��3W�-v0��A�y]{E�^!q�n�)Q 2�)��̖����b{n0U�[=��켿nط����ӱ��7s���O$�P"�e�f�I
ԦU������?�V)�����)���sN���`�L1"1ǭ���6G'��Nx��V'��@0���)�N�y?���ol�%+@�Ǹ��H�Y��å�<H��S;�rL�*�/���1�(�ZO_����0ţ?=��<���%�0������N!e��1A5=�Jx%�f�B�̸��A7���O�;9m���ӽ.LI���h<��I�^~o?f�A��;/�U��$�����}y�&g�-dB�=�2�@���>����ܺ;�p�B��Y�tל���(k���]@��������䦖z4a(I�S����x��p��L≣�w�=�)�x�'�(����%������/�Sm�YY�b�oT��8)���2NhȌ�L$�~���:	���@F9�.�h�� �R+�O�"�nR���r�?�d׺d\���p� @�)��-&ݺ�_*W��n^J��Jiˊ86��3\��Y���qr�A��)~��4��V�1����ϵu�8O�|��_mXƕ@�$���Hͯ6_Zۦ��!^BI�v�l�Y�%pѤǸ_?�_����nP��V�X�2J)��@�Y誏ʺL�ϝ쿖�lf��`�j|�+��9�Ǒ�jY�}�}�/2(w/�%a{��`�̵tØ��9\k���I�������H��I7��
kLu��-�,���!��{���a��@��n�U��V�=��
}Y�o�;o4T����V�k4ek�ba颚�,b�d�x������J�B'��+�e?c�1ā3E
$5�V��ME�g�[iN�,ũ��8_�T��c�"�
�T+G�y��W��Ɖ	sג�Z��w[����� Z��(@�nQ����1����l���V���x�xX�e���=qGM�ԋ������*� ��:�ت	IMl�$|Q~Kz��� t�t�&�
��:����˺�w,	+?c*2�l��	�)�.�!�1m���&�����u%�#7�f�ǹ�ب>)=�WK��S:K~�V����G�e�=2��.4�fM���p^�nS0j+E<�l(�����|% 7��g����CR�Q.vD&˓gn�Bb�|�h�A����d-h��*Frj_�)�
����ej�HC=�a��W�(�{�#Z���R'�8%�'Nqc�5�!�0,�x�����V�G�DnIX��^��U}�s��@������A;^������������o��Sc���oaSVb��U��(�	�](��s,�����}��H[�DUn�o�	߷:�t�G#��ZR��J��M�C��K)����i�l���;{����v.7�=L�y;��#(K��:�Z�qd�4d�X�2���ڄWXa�"7d ,P���9��V��#��@&�̓���I+:	NWҩ1���O�� �q�kk,'�_n����;hx@��Ӟl,��BK�!�q��g
g�n�8��$��:.VY1��"�lX�������^�n��6?A�����m�:FC
�.���޳���P�/·#���5|�����s�h����F��Z��O�CTY�m�<���.�uQ�@���\��MQM�TW)l��
���ϖy���	���궺� w�5�;�gB���b!H��a	-״ĭH���)��Ia@�	z��N=����+tƟ��� Y�7*Ƿ�J�.<�V���
����}EȥDľ��Wڵ&�0�2<uU��������.�J��p�i�W�,�1�������Y��u��Vѵ::b� �$�=Š~����}��`��n��?�dx�~������FpWc)-g-ZU����c�)�F �p�4O���Bs�؜V=��g�M�Þ�K"��4�#���d0�)���1�s��
�=�!��Y͏����t����^T�a�z3�b�[B��]�X�2�<�M� +vF)� 6z4���yqa��d	T"��\�npR�|})��6�o.$�޵�M(��yX5<�f����@ %1[%�Fġ?� ��m�C���|�7@S��vY��Qd%��UӲ�xқU���I���s�ϞA�۽�j��To�ta�K1��mH����\n�	e�DV(� �(.�A����'��8Y���"�'q��Ћ�$�t�λwΪԷ�C�������QC�j|b">p�+��^��oT���b\���#�u�R��Z���-�.cQ{����0�t�?��i��C{5��A�ힾ��bn��(!AK��6H�7 -��ˈ@Ӿ�1B�Y	CU�Ԛv|Vy�9�ӧӡP������o�O����Ъibל���3����v� }p�)RS���m���,μ2?�w��ǯ}�סH�^J[^9�yw��X� ʞ�6=������vX�t��Dz�f:e΂��[Ď�ɬc���0��W�r;sJ�\�����?�w�8��,vy�D����[�,�' 97v7'3��s�H�kY�yߏd0U*_�:�З2��;�+Df}�>�)R�_�N��SR&P�!<�� �s��!4nń��kT�C��y�Ҽ���ԤZ���?�*���!B@�Gh��L�,`�m��KE�0)K��S�{�����R�i���*A����ҖL�PrW�eJ/��>�a�5�{�b?���
l-O���JX+y���
F�:T,J.�t}췏[/�z�L!*��N��kW1t���-�<A-���-��I�И��(�+���õ@�s�[0]k��nV�)�g<��"��"i��ϡ�mrD$VFj��Z��~�hx|�Lv��ϴ��x��VV���F�:|Z`�rTDY������gT�q��ɇ뫦+\�)��l���t�
A�ݏ�9&���>�&"*���qX��0��\י�ߨ��,n����� A�j&��l�� ���g<�!"��}�`����h��,��"���"�4<�p$a£tJz����E�=�s��ŸOw��/;�;!���9�g���_+�����W�m|G��e��������,{�@(a�[�;�%�)�!�8�k(��b�Ac/H���i�x�T���-���.R
��L49,��Ҳ�ӶF�đ��(��i�>T
*��3��2�u0:�8T,&_��t��VĲ���A|*�yMԁ�q�?��	KQ]9~��#���HĦ�lV|�rXc�,1Ԁ�~\[r�ɘD��F��y���0)p��8Aͦ�1Q����ާ/���L��yByk�-ĸ���.��z4�)ǐ���s�|-���q ����n2�.D��6vY2�����!��/ј�vԒo䒹�V��l�
�!+vrM��y3���%�$u}vaB�6��h�	F|Ƀ�l
Gb�}h;�_橺�#ʅ�C��GıUREH���7���Q�B���_�EF#�?�Cs	��O�"���[�5	�=��������8J?��ȄT��q���w{���u�A7���xa��>1A~�S_"���K��#�d/'���d�/+f� s�hmc���1K��|�4|Ɣ���40���2��Gl:gG%�	�j�m�:��s_���(��/vDz6$K<���qr���~
�¼Kͱ[���An[�lx���ȶ[���2�� )9b�o�&�v��yW���a+k[���I����Ս���3s��m|�t�Set��gF9?�W�u���_�6UG�BS)t]R���r(c�֣:��@����!j�":�[��M���1j8�nh��[���9���,�����AP=�7ډC�v�B!��8����63"%OoK��S0�u�6ׄ���ʞ�^�uRB,!�ʊ2Z��vBơ�7jj�\��Rj��.��*6������c^�%��K�
���F4����~�9V���RޏQ���b)<]�u�°OJET�[A�`aJ�/�n����8����-6���5ƃ�X��ze�m)<p��F�H�
!W/r=4�SE$Q�]�i}�ɘ���m����0¤��_��&/��o�׻��A�Bf� �C?�KtM�X�*���>�r�+�D�8!vp�nWk�]eȼ:�FWۼ��V�=!ӗ�^��R	C��/כ�.h��T���g��^9��7͠R8��i�	h����;(���������qc>Δ��Cp?���eД���52�\@c�@$����G�1�J>�Žp�4�.�}�c�g,Ԗl[���{�G��U�ꡫ`p��Io�~�Px�n�qH�83i�"+m�(,�C,����1���~+��yG�M��%}�>�3��k�F�v��E��\�w}��Z�SYg���B#��#�-je�"��u�R��g7B˞��s�=e�a=�#Q>�}�0�7�qP�'	<��G��O�A�oO�>NX�G�CpflF�[׃}Q�|���KC{=H��������|
흤R _����3{�f������#�R��Ih:��F��Oϱ��n�RE`�&Ak͐Њr+��ǍPGj�f �U^���v�YZ����K=�eI@Z]�ژt���/-d�����XdxV�{�h�Jk��W�L�oF�WAZ�9�-��"��S�Ξowx?��\;x@Jh!3Z|�'d&��?6;���B@���T��i;�X�s6Qt�
I� ����bs_�OD",��<���E��4�C������G���hb���iK�� E�s�=�m�S��C�E���/r���<�W�:$�*k��s�Npne����NV��r��\k M�\7�0p[�Pˠ���
=����+�t�0���$�G+ik �KYܠt&m4~�9�Ot�ôT����/�c��c*h�w�<�$]�3e2^�c���wx���N�cI�ƭi�\�$&��ޟ��<E�Z��Ebِ�oI�i��m�gL��|��jV�MۧZ DP.S?:�����Z�����G����)���	%�'5�KS�j�J�-p�����L�h���P@�s,2���S���,%��zA��-�iX �
'��;�Q������uod8n7n��-�zX]�,����
��)���'I�lv�.햶R$� ���-���7�*����ƞQL3��#Lz'��Y�\7q1��g�P`�u �W�g�_�p�&)1�D �_7k;��8q/K�>]*��
#�O"�n��#8��fD5�U'O:��_xa����x;��X�Ig��Ào�Y3z��it
�}�R��Y�OL.v���(�syn��$�.TH�~*A��3����vhU�N��U�:C���O�L�Wv*��,�z咠�m��ׁ��dӞw�h�1>w9a��M��������ڋ@wJ#�͸T%(�c�f�t�*�Pjs�7:���ׁT����Ve��z��s������)�s�wd�X��l�,��5G�ǴfL�*]��E�7a#�Ƥq��5�C��H�s�p�
�/DHJ����T�y���۾��^(z�UGnd�cs)`�̫��h­S���h�[ɞj�j�"��ZX�$o���ˏ#�a�c$X��G6ɖmv���B��%��:��)W򥦹��SN�,B��vv�ǆ�t��߮�}!�J�yd�?!�'P�[�<�WrU��S�Z��9��!lߕ0Xלvg��9�T.7Nm��t/�4w6K�N���59&��],Í��bv�HU����W�s9�񮬙�����2D:\�b!@u�WmR�K;��ٛ����hDMD1����<�.��άF�Q�u��<�?�s�V �A�y?���: f����Uր�c�i�"�]���J�TɂǙ�n+�XC�����#����BL1)(A�J�Xd\ͺ����ѯQ����A�B�1���	D-i�p�Zj�j��; Y��V�&厞4����&;)�U)*���m1`ե� �zB��cs/�oΌ�
�J�'U
�4��B��^�y��>�C���)���17���P>\�{��r���r��(:���.��q��c&1sQm�C�[���Q��:���,,�4���~BEtZd���(pL�ߖssI�!��!F�`˂�m!�����vѨo���=��n�׍�1�W�|B��5yQW�������nͅ~�=^�'�#��b���y}��v��&�G���o���a���W�*$wݞ"��|��y�m$�
qwߟ���|��e���#_�+���$�EN��?�N�{��y����k9q����:���Qgdܫ���BE���Ա�+Q^�D:X����4��9}>���Ʉ1ه�v��a���lo䍾��&3�k�M���!o�3�k[2Q��{wp<=��Ц�YٌE�m�l�]!��򁐏U�ng�$��u�^�m7�>�l�R���n�V]J�[c$T�r�9[�TN�5w4�᧑��·�}�F">`�k����	�0K�R/�	+�z$��6�q�H$��e����#x�j��W��[ ���W�3^>�l�`�fV�������e��0��Q�+ހ,����s�e�֒���D-L�I#cPA�S 5�q?�$�pBf�򐛠s�G�g�>:g�6{rR��I��m����]+��a?;-%&x`�W��y�1A�.g��Ul���ڣ��gs��)���:�nJ샥&`:����������}҇�����q����Wf�.r�%���\�ѷ�ML{�\>�/g~�6�I5-����.�p���� �7�h���w��c����j�yH��kE5�S�A�\~��o5k��դ��)3�����n����m�UX�.�<��&�����EW_VPD��fFW��
��,������6}�:��L�A9w�s�iE��߁=ذ:S	S��̭�F�6
m�:OKLY�{�ء�v�,�n��$a�x�F		��ߟF勮C4QR#��^��=}���+���m��7�`�;��E#�����SNh�_G��@��� �썯�	 �?7Uq��f�
 �4LEcQb|Br"���x�>U	�yܮ�H
������_�l<�k�}��f�.n�:�	����e�ѫ����_frX.<Bܕ�KQ����S�pZj���3G���iȼ�G��,���D�.�D�Y��!��t,p����������W�9�4��C ����;����D69p`�.� z_�4J�M�5C�x�'ԈӘ�]�>K*���ZD}*w�֒o�(4��1��Y�am������k��.�I^�H�&nf�݈2��N+���,~n-��iֹP�7T�6����|�Y�0^�A����NQ�\&�u�B�to�V� 
�/���Yp�g�Ȑ�c�l$	�x������B>�������z'���N[�:yg�T2ٗV���r(ڹb1�7��43V�ө���|'E�oK+ɏ�c��Tг')Ә��E���kt_�3Z�8S��u^�w�TX��g��ȾA����As���[.�R�n4io[a���v�YH��ޘf:7.�|L�<�4�ע��������K�~��dVNj�X�)Hђ�n��LՐ��w`)>@�<�T�:��\�/���qZD^�OMe����z1?�}��R���f���=��w`;�u*= O����Z�pE� �RwѺi�qDk��l����|P�@�u~�y�������rItw��|���2~�Y��4L�2Z:pt��#Im�9&ԯ�C������a�K����fgq.���{Y�=7c�U��{��ɓ|��5�����o�,,��P �4�w'->$��3�w�}�bߩ���2k�f�Vw�ʄ��@֌���*�n���th�X�,���yV�#� 4c��yS�.��~70h�$�_p�d�{#zˁ�Z0�H���%?slF]|��J�ol��(���1d��Z3b�Dm_�vǠ�d��d�hk�8u@����(��3��8�訛��e�j/���z�
&�MT�l��
>���.yP�L1_��Q_�x��?��FB(���8D��s�����Q�o-��0�BOH��x�ow��lv�G@�S�)����#=	�
gr	�y�IgE�l5���A��fD���퍸jh��X�^Z9!.ē^|C��-�|o��{be��$��xX:Je�L���eYpY���Z�覿�uh[�(�^#Si�y&n|A�ih��z'�0��E�e����ȷ�ʟ��!~�����Ga�{V]�)�����b�B�78f��K�{���nqNϊ�";u�y�"��F)���{���n��ҽe���!����n�y�Ct�LHwj;��`����r���������br�w�c�6Z�Ģ,�LD�G�V�w����b�i.��'P��Y�%�1R�)C�����<��
�i���(����Ih����^�`c�1	^6�Pƴ��{X@��K_���
r�	�C��
´:�1Ⱦ��D��\��\�)m�������<��:�
tp�Z7gl_y�gh��N��2q{5�vfYF�����۷�d�{������z�_M3�A�U@�2˩GorI
����	
����B��Od��;�Tޟ#����YOq��j����2�խh�[�-q�C�S����G;��EC�m?�0�̐b�� ���kf��.��>�s|��7�����hK�s��͢|u������3x�z>$�������PK�7fK�h��WZ�[��ٙ��("�BC�@�<�@�!UK�hEj(��Ѳ�j6�/����n'�!O�#����D�=�am�����[��N\��I�G�x)�|܀���E�,��[��S�dV�5�j���ۢ�l)DW��FĻ�:�sm(�֪6�p+ef\4h}�_M`v�B���<��f�B��GP�Z+8~}�?j���a[��Xȟ<��QV%��p�6V���k�&tj=�P���C��,ߎh�ë����}���yK��.�9/�V���,�:_���tl���Lf���B[:D'}�}صS��֛�cc���p�z"��<WUb������cN+hs�?�198�J_;�uF0�l(�ޜ��X�T+x�[T>B��PO����hTe��
-t�`��)']wKc�O6�19�a�u�,�uߍ�KD�V���St�*�k�/.�g�j�(Vs���R@��O6(�c��V�Eq�:Z�TY�H��������N�6�h�ѣTL��é��{s����	zu��=c23�c��h��C觜�o֒!�X�^c�b��L��Qfv�����ة����.�%���E�D~��]���a�$2��kΠ�,)�_T"����{QY�B�a���>��cN�K�@3��(�UF��o��ר��8M
1g 4u�~b��_��Q��E
-�o#��	��$��zԜ�$՚���%��_xoE1�����C�CM(��n|X����$9IN�i[2�~
��4L($�i���z�����X�9&���C 5<���Rũ�gD��Q�ֺ0��H;m�
~Vg�Ǘ��S��Q, ��I5���K�p�RR	%->�C�V��ݏ���^L���?�}� ����Y�d�"�`�rZ�z8�{{��W|ũ�����p�C��y�&�Z��2*�{C�co�M6������?�Цݛ��n+�=�E:(Vls�v�K��Z�Yp�7�ҩ,&µ!)}V�X�-��QN�F|���#߅�Ώ	5/Z=��5�M[��)#Z���얷S��U��LZ�ot�0X�<�u�9�ڪ�&f�~O��e��냢M�8)�]F�t�25)MP���_��x�p������	����A8г$�f�8�l���`u�B�5��k��My�����������XQ�� ����A@�F��d�ƶ��x�E�z)R	|����=`<������[��/ �9J�<�4���?�-��ף'Ϧ�޾�gl�S��y!���
��-F�=�Dk`���\+�h��}*�G�g�=�<��]�Gl��]�q�r�l�
P�y�b�=�J�t���4�?CNB)#��X�G������2�u�B�+j��'�q�l��:*gͺ���)�[�Cϵ[���"�-�{����	�p����_3�]9��,�d��7<X���ĕ9K���Y�G;��7�R��p���r�0�/�KD�S���ߘ 7̃X��9�j^���ȿ�u|�;�q2m.�y�*�wuL�uB�M��	R1 j/�
� �F5-ɿ����w&"Q�\9͉蚍6G-F8t�@��D>��)��_��w�nNc-Z�g��>�D�	��"�~NXι��у���U���	�K�����1��ꭖ��I��0~Ćd�r��3���q���$���쒟����>�&	r]� �J֫�\$䠉Q��] �'���� �qTb�i��.X����i�;����^z�<*\)Wl�FL��>շ8P��� P¹���a�����23Q�R�l�����`�oHGr�Z�.2��i�bU�mfm�dq�"�6���`�j����v]J%�6�!3�y!i�.�E�z���z�����|�3�ţ ӖM�+}8��M
�?��� � p�=�*���u�M`F� �7���k� ��p�'N�T(��{��������eͮ���(�.@@�;�q`�51��̇f�k^�ȭR�sR9����e�c�xw��3��������U��ԭ�?,V��`g�m���E��fװ�����3�b�$�� �H�!?66�:=���ݮ�f5mgm��ej���"��ƈY~�4�M��{߱��N��@���餠9{Xm�(<�e�b�������)I��)�[/�[��̑x����T��m@V9 ~&9>�F��f]j�*�6l�$�i�T\!w�B_�c�l������j��!S��v�/ʳ�D�-���ꥁԠ���2%�-
��{��Dkw(-d7���N��?Y#�m�W6p�q�)�(�̦�x���`kufh/���7�����j6Q׿�+��8Fk�t+��AU�g�N	ٌW�3�Y������G�B &�&�ށO�ם��u�C�a���z���ug���ɞM@�ܭ�_]I����������o�,�����I6��+Ԕ��r+e��w���j&�_GJ��&i�Z<_2]"��G$�k�M�)��h�N[��_c]	��������fl���чNj�g}:ac�����,�l艭��7�M	�M@�u�8[��qQ����^`���'�X~G�/u�D&�5�[wg5��fMPh�D�C��z�,q2&p8"�A&�]y ��a��A�s��w����Nv
wVpI�t2y�p��j�G4}�{�-rV���x�
Vg;|P��8�N�y���� E��=��>��:�B<�n��t�1�n�{�:0��\^�z2iq���ԭ�P���21�svG���*�7�5�t��p�w%�<�
�mQ�Ő�!)���:�P�Fd	4�i҇��-��=&�t�p�q�E��QM�6������'6�<s��<���w�F֚��C=���,5	�Wr����=�
V;���6"l*p���$[)gs��0F��po����(,~$��q0���"�!/����?���<��W��7.�`��b�� +>̄�B�t�I	P��G&7Ä-ƖX�=�O���-A�O�M�ʟ�Mo��C�����e�G�GP� Sv7a������_��yﺺm1�j�����3���c*�M�k.)@�1j��Z���m09�G�n�/Y���q����ӹ%��y@=�$�2�T�X��{���/r:��ߕ���#��H��-���r4���H��:	�d)�M:�p@W�\9|�E���ٖ� �ڗh��&
���1kc�%}D:�y���D}��oR���$�9!G��
��eAk+��6�DA�P�F_9��j�A]���%�W�3w���s�����J�a��Uˀ�E>TjM콆}�=�vn�."�\��)6u�|��8J�.���o�?D�`��+��s��������M�.��߫������-�9�q�_�*�m�W���u�D�G�ɶ|d8���	���ڝ\8��uSlVꅐ	!�lK��`W+��cz��[�!�#�ϼj��,��z�p��WM�8�԰���
$w)Ŧ�:�I0/L|[��m7W�}�hW�.҉�DzL؄%���e��C��D�e����x�E|\l�
�a��~�-��Jcخ���SfG]�Q�sQA��z=��$D�i��y���p1�=~im�ڊx���[4�l�c��	�I|�) ��
��&�Ϭ�C���j a�s+J��л�]�O6��LH��o�@��8*����,������]�%�cAE�g��41��� {�dT{�\� ���jG�S:c��O�tP=�k�x�s��o�&�J����NZ�A ӈc_�]�~�٠�����R0C�B1�N9�V��+��~�9f�j��,2Z�_�"�����U�\�\�~8�^n�h ��Z������P��󨁬{P�k=��F�4�9���c��Rl	T ݄v��\DE	"�vz��^��:ؼ�5BL�=�]��M9R�w�Z^�������F�K�����b�z��Ӑb� h���mܢr���?��/؁o���z�~���(���S�)���� V��Z�����!���~V؂=<���+��Y�I�#cP��g3�@$k@��A��K�F�M�%�"�?�Z<11��G��� Y"k��P�F�C��b�����L��39$[E�L�Y�!3/���*L���ʺ�z�1�{םC���D��f�Ylמ���L�p;w�ˎfL�>vE����ϭ2�r#�`AKW�G�RƐ��UyB�\�j+<���,�m#��*w��=�0<�������<p�\�#�Ti,��6՛a�g
L�Ԅ�h�7�jE/yb�̋GeAxEjF�l]�ᶆ/��l��3�4���<)<�CksQ��̧���>���2!��Z�Y`���$�R�k�Y������B˛����r����hЪv3��4��[\O}�q�D�i�b��Z�/%��M��۹Q[(��l8yի�9���0C�Lϲ��,$9�c��%?41鱪�ĸt��T��S��ڟ�O���l�Z,	X˾�|����(s��ϵ��+<��o��&s�6�C�~kY����w�Az�.z��xw�}��5��qc���
�h��7*�skxe[S�	M�Òf�s0���M��a}��%�Ҙ�D��Y��{'d�|�kw�P6�\���p�G]w�q� ��F�Y a�H̄��wk�0<�4}�v�o���7�Z_�~��0��{�}��?9���Q^k ��e����G~r���tK7w�0�aw1�J��0o���@ۣ���2�}�6@�?i�5��������&��o�I�Ĭ�;�H/�3i��z�V��M�D�I�y�I��7IA��<�x�-p0OCX~�_Q��Yi��V�=��[�jd��˒��t;�7�!dkd�#���	 �!��h_)<ޏXՁ���L�\�F�CV^�)�����B=���(�1���Α�@J�ȺJ�p��g�1B_!vBa��>��Ļ�X���z�����.�&<����^���ZzW�ca�Q�VRC�az#�ۋ�R�lFPJ�8�_y�߀6�r�W,O�H�s���od��R��E��au"��������8�&#�\Nk�D���S��'e�]t���|�y)�O�:;k�cpK�W=~Rs��v��}�$،N!4G0�3"0�)b�9f�Ƞ��p� ?���?����BS���Ŀq���?����^-����I�
�2#�JY�u�#�{�8�M�ہJ����<$�FQ�%�IX�ʠ�W���KO��v��:�B�o��3,��7b�ӿVְ�����g�F���6�<��&����X0%���UHÿi��w9�c�$,iSK~sh14�SF.t>҂��w�v�ǏW��2_�;��bc���޴-'�o��+A��ֺp�@��GҀ�$ǈb?�J�����H�a���EM��e�d�/�X�o���Ι��z�O��wǩ�*��rj��>uJ#����!�a\�����#Ĩ,܁��!�C���?d�0d�H��͆;��*"�0�ٞ7u�]��Q�^o��ZH"��|QT��Ҝ';�"wmK|3���9�D̏���Ugma!V��!y��Y8��!�o�v}Q}��n��Bb���ś��o�5�D�-�
J���ŗ*����{*k���E8��i� ��z�α��G5,QH���ա�Eo�J��c��t>�+���ц�;��Arm��	��Щ�|E�rK1���Ll3F(���?k$�XXF���B_t��&��'���\���"��� �Kz a�ٌL����Y�_�ϼN/?��g�EjA�m'�
�3~é`����o$A� i����\�n�Wq�}�>\��I��i/ _��-�/yE++��|���$ɡ_��/�ѓJ�r��.E�!p��|��"�XU�V2�@Oy��	��ɌX�����b0H��r3K���1�z��ׁ�IC#zM߷�5'[��k��Ŭ>���4ڝ,;4JـN����d���q�����- R��C��@X��[??O��5���i��$־X�H�8�T�Ȧ���lj-<�]ՙB�`=m��o�%�
���eT��DȽ������O�����W'��̵�vƸ*�b��.�Ĭ/"���~��!�n�����Ǧ1ņ���vP5s�;�� ��C���/�z��cE�#�{1�Z�.�aI�J���m�.8Re� ���n	.�H6���� �d��5	6��w���Qfg�c�>�X���!'��	Q�/9�^5#���2��w��+xB��LדpE�-I��֧&,o�y�.:B���ٜ ܘ��q�FR�"�V-d)qUג�U
�8���4�7�\�"pJm+Ô�.g���o�"R���!�7��.�f�n{�u��cb��/�����'N���{�P���'�*7a��������A�i�� ��;r�C�P�PgQ���$f�n�FI���ܝK�y����Sd_�)bU�t͜hy���-@�h�_�7R�*5�j�H�u6��V�˴h�}z*'c�tka�4O��������wzqi��P6A^�\6%S⌢�h�n�����ReZ����������dy�{&ޒ��������y �M�3�"���{=+bD�HƫF;'����Ҙ_5�q�Ԓ/�PM�1�յ"�hNi�=��X��{d�a��3N��)�[=,;h�⸠�J��є"y��軶��@dK�Q#��~	�s=?�܇"�ͯ(2�ɕ�}�gd�}�j��O���)�������������4,F>�í�m���e̦
$DD�nr�zL�M�k��h*�z=�?��]��ͥH!q�E{`�q�-�_K�D^��B�Vw=�a�P��Z����<��k�%A�W�I϶������b��w�3�3��r�X��n��Q��0�`��Ae��k�dS����JY�D�m��Vp�$�!0qϮ��_�{��˕�x�s���e�{Z���)i�y�z�:�'����@���,�>-ѫ�aR�t�i�5룩�=]��1
�
2�W�/��6��ގ[{�����N"=�К'6t��ۣtG�P�ND󺫺�27��D;�X�)3���&��Y@�&¹%�eh̥)��$�W,ߕ��EK8� �;��۹��lH^2����'� �S�ѷ�4��/#���KC\t�h`�a�$�X2�()w�K��|�)ӻ� �g��n%�+�1�b�.�8L�wa�����%O����%j����>j�u�V�1�l��ߠ��.X��Gͧ~�Ŕ�6HZ�H�w�U���B�`��2�JB�S7c��]����8)�9ȝ�2[p�%��5^!"y!d�Dg=���302%�Zy}��Yz�e�d��9Ei�v�9��_˫��4R�P�[ �S�S����R6�Q���������\�A���M�_��hY�[�Gi-۩��膾�XLඋ�O���S��f�3�7�k��	��o&� \�BfO����� ��~%3��ض�
Ms;@C�m/]=��+��3�ڶ���uJ�s��W���3�*�b'�� D�t�;��/�8z�@2WWZ���H��W��0@9]5��C��jPrX� �8�.�1��W�_C�J�J]�	�Z�)�/��+�bT�[��,��43�s�ݫ��wBP��藦���Ѩ�����yܦ{:pPV���YY�jCI�~}m�ri��Z�r�E��C��4�`�Ьp��9��ڟ��+Z����ŏJF�iN�
���6@BN�s�w�؇�Q���0ÌωM^*�ҿ����]y�v<ꅙ����vY�<h�b�|��-P]D��B8�KO%�U#CT@�u��m�`�\E�����}�)A��>#G@/W�@U�i&�'U&�3-�:����ڋT���o򹦕�����o%��������)ԀV����(�G��k�TP�g�HK3�A�p8G6�?�=��WN�Y��K����u/	��{u{L��?byw+TX��pW.��9N�/��G0�/�U���bt�d�Cg`IrW����`�7�(�*��!s�}�����s Bߦ�|�w�~����S*=�9ㇷ��s\;+���d���]!�%r�kڽƄń�X����hy���~]�w���!�y������٤����<'��e��fO㎚�U�kE뾧j��4��e:hX~�j��И�N�G/�!̱�e���Q�R���c}�N��}�@ϰ̈́�-T#����^��KTzG�y��[�v�1;9p���  ��$|�`\�Z��?����z#�^�5BCA�#*�G�.rl�T��!b+N@��}�I[��6C#���lW�Ǎ�y���9*	�>��Y/���K�S�W�f�\*�=k8d�o��)���O�y2\��9�P3*�QZ�������B�B��R��]φ���&YM�ﴁ�O�q0���QmB��B'�Nu?G��%:�_�k��x�q�԰VI+�p�BG&*m�M��i� ��h�F�t��.�����BB�-��$j�uR���F�pZ�R���ƈs�?k��(�����a߯%\�-M�B
i�t9�۬����R� �_\lH�������&�ͧ��͊h`���Ǜ&���H2��0PL�)NH�c��I"��.aC�G�U�o/�\�� ��"�ф7����9v�Dh����������v!V1� �y$����ٍ�[����}�F�%p:�1����;�� ������`�6fN�Λ���R�W�  �̖�8��B�<��y�E����f�����P��(�Aj��D�\�������cH��z�{֒� �u���/Ri�s�k�����`x�%>��֔(*�c0������72�]Q�2�td�H��j��'L�H���)�-Pj�O��/J�)����|��c�����8��h\T�M�u�������F�[��v��E.���>"dy�nP�~}����?�1݃ۡ����/���\��xgyLI�.�*IҴ]���6i}^s�gԞ�Ul�������xM��b�ZD��>������q��z�K�Z(˝�����������Pq������6�n��/��ށ�ǳl6^�s��X�Ӓ���}���7�E�����u���猪]���(�мI<�c�ЉK�P,#h�bY$y��������n���V1�^nc��Kx{V��'����;4�<ic ��}����x� @����l�I���jݯg!�!�,�鬻���v��`Eb>�B� ��~U3H2Y�1cF�|P_�mui�{�����hBP�u�)�~G��Ey���3h>;ف(u�	�?4nx��JRt���#[
	��W�3�.�\��&Q��{���A9בW�o��w��W�lX9Dk?ә���#��9�����J������*�K�qY�	r��m)�#�P�7�/�;Ì'�b'�ݾ�*g��pL}L��9P�ꀴ4DR��)��Ɂ+�SA����凱ͻr=�R?�B ��!'�6!bߌ��}(��5B��E����#h�� X���S�R��y�:�
��S���Bg�� ��{�K ��Azp���ߦ�T�=&�J�t!	��1Β��%/x���O_�~���St2b�-�I?Ʈ�J&�8� �20$$$�8#�M~�$Ofo��)�����gv�~���e.�:񱒉��6�LA0�����h0'/�ǾyP
�7���v?��Z��Qn��ۯI���_J��0��y�u1C��B��@y�h��{�!?+R1Z�řv�p�A�)�V�������K��L[˺�x��8��9Z��.(�9È��웢�S]p+];?�jD�׏}o��fL�wR�M/.�p�E����D!�j�;�?9N�m����2_b���4x�?�0�!��ߥ5�/���eTυv��B��s�!]Ҍj�tDf�����ֈ%���d��a� 4Ђ�tH�pe��ێq|B�{+��G����cU��ɔ�/�O#���O?j�n��rH�.W��.�T���4] ��|s{��N���͍3�$2�:��������C]��L��y~7�_����&�$���t��0�F�||,G��M�]�K�9���_5��n/ڽd'��3
�� 2�ݠ9�	�4 0C>d��5mj���+�ݸ;z����!���nZҀ��-��p�_|��{��N+��Kr��s�AYX��i��}��U�"g�QSUH�m���%�ZNJ��A$�Y�	�Ф���5dQ.J<�X���e���s�?�m\D [K�����^�/VI� ��]����^��R��i�!7FU�݂Ə�_nƹ O��Rdц2�U�S�5C��XF^����/�=_�;Ԭ�H�kGC���Цf��cX��4�wyY�j^ˀNTCV�m�D���N�����be|n���kG����Z�0&E~^FSw.�h-xv���n���#���%���4L�P����D�� ��k��Z]�~6�i�������e<�[���G&Lf�����lx5 f�.l���SF�r��h�N���u���m�	�W���CN�:C WL6�.�����Y�$�y�\�̵W�je7��H
�#��|��8m���/��f3����S;�C�>��9���SD���a~�Y!�v(Q�5�)_�����b1�}Kn_?����\שj�
���Ѓ:���9�)�A�[i]J�O9LEw .�<�~~
�ߌ"����K\]��N�W���%NZ-�؆�7���mlm`)|;��r�N}�+Z�=�D4��(��A��WG/O�?���w�[?�'�)Bb��B%v����ڼȶ�H��(���X��"p��/������$��EF���!��g*Ɩ�"S`�y�ۉ����u�5f������9��
��F?L�>	�Ӳ��5�ʁP�^�$��u���hB�8[�/:h�v5l�5��
c�S	���g��
�wM���d/7���,�����'CPϢ���<1��������D���9Gi/1�"`�o��f�7+�K�~���;&��b3r�T[�d�g4���]3M�uE\%+�o�

���Bv&K�=#u߱WCg���nF�o 徕6��\��[�JS�D����P���G���Rlu5Q�(����6v��^�jA��X��k��[���R�c=�_��|Z��þ�f�
�ΡƉ�#q)��4ӗ���ެ�з3���X�24���K�
d(���Q���*�1�{O�e���9��j��Y�|���e���;{�ҺG>3濸��+,�T���a��J�-Y�5��.Q��v��ښ
����xK�_�`�&�zۍ�u
�@SN���V�9c�< ��/����RR��K%���c����;=<N#ȿlx���q�Մ_+x'��;�'ȵ*����a�z"�[C���BxY-8s82��Մ�h������97�Z$����E;t�Z\E@T%��Sh�EDcD7C����K�E��2)�H�8,��R����6�7��!�{ĥ�l$�-� kV�+�� LI��
�9�K`B�J��/��G���
��F��B2n4�b%>ϝ�^�Q�Q�Co+���5.xӆ�!���y��虗q����ojxU	S�Q1'N1J%�ZU}ħ�v�n`��I=G��Lhi��OS�u�s*W�}$q F�Hd�^j{�|�1��U�a�o!��!�b��7����ae� 7o�̇B�+�	Vڠ�b~�)��>���tMh �0b?KٓXW�p���qrb�j+l��Ԫ��[#��hh�"$�B�z�&S�m�T������U�&�fʇ������VA[�cR �V���#��K�9ڪ���W=����{U���[%.!�!����!�~ b��-��fHWt��Be�r�,��,���'��%[-pQ�N���$��%=���A�Q�k�zΆJǛ�)N������Y}�w�_��3�
5�Ax��+���ȚY,������uc�дw��k�l)i͜4� �.O�=�W������c"G�`��DI�����t>4AN��Co.��B�~�;v#�V4�F�ny��R�v Q>�<���I2�����칟Z��CQ<�� �{(.�2��O��3�#\&��{2�~����.�V��6������b4��|��#W>Y�I����蝄�PJ�	�sQ��F��PT2���x��S���F�q��V���	�G�Ny
x+���Q��������瀞��m�n��^ʃ�$�$o�Hj�$�N�:�`��s��z@�����	/	���	�~]7�uVCd�A��x�T�%����/���|[�N!�Yg/�6W�ԉ�΋�YL����G���ZE�.��q��`�A��ux�����J/�my�q�!e\D/5zZ��mU����F8��G!TSڬ����H�>��4��8 ۅmů���V�>A����+��?�(�߬�nj��b���L��*�"�s.�:�� 1U!�m8����2�CQ�Ae�B�Ihҗl�p%�ﱡ���ٶ��vdpl�������#.ǫi<#�:r4��\;�h���,q���� �Y�~�S�H�V߰��-����7�QG ���rop�Đ�`�P���w�eg�ZB S��:���=��H |���H�PL,��3��[ae"�d��ۊ_��c���S��A�t|9(���y
^��y������/����P"����ɂ��nE�\[�N
���KnC6�V́4���NM5R�@�
�=S+1@�RZ�H�S<��^���鱇���'ru ���v�S���!g.���V�TK97�Po�n�>1Y�M�X��a�=Qݮ���B���?��Jq�p�xS.���'r���O<XXf��/	T�wWD��-�1�J#Q3I#)��9���Z���_�+���bn�H��E��8�<q����&#	�����6��-��H��~��9�C���b}g��PG�B'9'���咓����e~R����ϰ�*��D���it����`�ǫ1`"
��П;�8��➴��6��*Y~kx���SH�BwgL�	O}�$A�8=<��X���=��,��6��"����5?Zx�V+x��S�0D*; ��-��������)J��_���ƠШ*Js����
OU;�L-�ngq67;�:��v��Š	�!�/&G(i.xQ��F]u����Im����մEI��#$.)�1J����A15�'��Mc�6i����~
������N�J���,^��Պ�u� �24ZkG�dzNd}bͷ������@�7�`c��F�p�|4V!����\f��V�JЁg�$U�=OK�AOR�)�SÖ́���*6-������')���)���&�q����^�������l��H?�w����:�ʹ�����w0�(��+�)
�'�zE('�ڔV�f�2��3r��к6�߸}�Ǉ�����;�zhD ~%�l�Ȣ�E����*o{&���̋�Ԡ� �&f,A���:���3e��w�E�k�>���9�8I&\���T��oS��S����s���#j�Ak/*�#��$��x�ɠ�{F��򐗹͝�c-+��Kȍ�����}�K�j��ZH}a�ϑ�� -�	��Ձ�C��hc�o_
��ߌ���눾�D/�L�RehV���j(Ez��Q�(p��a��Q)�*X`��2<4_�=!6�.9Jհ��b���N*��l{�v�\.,;����|S�X�fv�O`H�Ul��y$�!��=j�\$��]M��1;(��S7;PU�
y�ۣ�3{����1[��cd��~�:�Y��R���g�M�1'���gn�7]To�T��b��`���Hr�C�kK��>�3�}��{X�i5Oع��B���o�������B|I��Jcb���C�9�|�O�ҥ�����$�ka��2�0���Z�?�:��3��:�����I��)��yeeSh��H��b�c��~s�,)
zK��ld^>�oE�@q�Qh�/�(1��:�0�NGES��r:��,�fg26�]��OO�O�� g&;�`#�-��i��]��x����@k�f����W;?��|L�RX�Ѵf[�ݽ��rA������r�Fk��ۂ~ڸM�F��X��C��d�%-%ΰu�p67Jm�6�˩{���t��:����G Bf5jF��`��	���1�]6�^tc�↥�Ą"h�j���m�j��P� -��q����[��c5�dyh��x���ޠ��I C�\Yþ#�� �;����baA�%%��d��NӤ��3t�iH_v����U��Bt.�V���w����Y.���g?�ЅǼ}����j���1�E��S-�AT?=Z���V�~�3�{�f���E6��pp�<6pAk��������.�Z�PW����g;�l�h���������/��>ht�8^�n'�� o�L�7ŋ�c�R�� A[q*���K��-U����w�FXܓ�V]�t��̕������}#��-�]��;-����	��D�d��d�l1�m�J�|uE��g�.�͘ܧ��s��|r�����W��ٓ2GWJ̙�U9�!Rj���v����;�	�"��D�evpP�x��زʵ7��|+t�/�+�~M��
��E�!
H�;�x��(��d�����S>�~�oɥ�ź��N���tĒ��ݥ�<
�0�F�'32��
_n��j�����}_"��n�������� �ѱ�T��*ۡ[���a��4�OF^C�g\��i�q���ܔ�f:�[LX	 �z�u�X5�ڟ� ���+m>Вg*�!�8�!y�B��?�X��8�>�K�	������?o~Đ	d��� zŹ`0t��*kh��`�A�^���z� p���;�3��^I�^L���`0d 6#�ۃT겾Q�@`��"�$-޽A/7�jy=(�ؑr���������^v�9" p[M�����D��V�P-DQf��L�h�$�ܭ����g��5*
�t��y��ƼeU�و�������5�������υ�Lz%��"ҩ1ᨪ���OɽR���E�~����nɾ-�]�/r�p�-E'�o�
�2���(t,�'����P�BɬQl16)8�/T ������թ[��s_�A������!�q��`Tp���XWOn�O�އ��Z�ő��kr;��v���^k§��׼#[u���ǵ?P���ϩ
��7F����>Z�O�f�^g��-f��n�*L� �)��S�B0�%�W|�C�z=���C@V�1l��7�2/}RIa��1ع7�������Fx+ /�K���挍?���u�@�}'��d�;9����,O<ȹ�B}�n�����K�O�#@t�c1��L5�񛞠�Ȥ5]\C.�ӜN��G{��ِS�IMvvt8��}�ێ���EfZ��Y��,T
$�ؓV9Ϝ�����=�;�sXB�0R.4ejawz�i�g���8J�^D �T/�_i�l�ֻ�]�maw4Y^��RH#��vCg@��X�����A@l�P�t֐��#�1@�F�p��2���>FK5J	�z�ه�J� ���ˈo.bķS$f�J'H�j��=�F^���t���Ul�lZ��ґ`x\��d�F��ZD��h��d������3cz�.^���5��7�oL5eI:�gJ݂��CZ_X�Z�4����<���*f7 	�V�~���h �[Y���G�&���׾u|D4���s��H�t����"��K�������|0�5K��2��|�T�,|���f�e�6�T.v\}T7�S�W`�iE�X��gx�����3Q�Wm&�<;ڧ���5���'ŏ>+�
��!Ɉ�Uu��!LS�&��ٟ���d��!87�Xr�C`j���T�b�O����M7�Ud�	VFI�+R���Ka�D�h� �F9�.�����+7�JF�e�pi�e<�G�HW��ʙ��s*Q����W�!�4M�~��ݐ<(��":C�w��0�x%~�D5����/#�Z�rp��;��V�dA�`W�h:��e�H.WQ��MW��ں4\޿[�W�\�g b�Z�v��.�a�c$j����X� G��\$w�N�5�wK��m���M�^.4��zB�@����A�65"���[��A���ľ��o���;,F�����jeQ��h�T�56_o�=�D&��l"�{3�st��b'n�-��.��;��I�6_J�TUI}�6~���vނCՇ6��
*�5��}�46Ue�ͱ.�${�c$Q
n��.�7;�n11�d�,�@�ה?�^5��זjh~�E��ID�n�!��G��^����\�g�< �p���D?!�R���;�����s�����V�N��z�R�����b��Ɵ�)�ʻ�BC��jI�;y󑸖k���X3*����Ѫ��7%���r���(���:*���Z�$u�DxZ|�*o�I8F)r� P6oU�N[�,ψ�{�eޟ�)� �jC���L���%$��tz�{�/d'�>o^H�˼ �yF�`�L�Nր�@�+�hp��ȶ-�U 4�����N*4O��`5�����P�� 볂Pd�#|#Vk~�U����s|�� �㵯#]K�]p1�`�͛^��q�EW�֛Ò����Ѥ(a�H,.�ɥ4yj���2\�h�,k1tS��R̥���O�����8�^���~��h�oIz'���b���f}�Hͅb�E��������y�|r�L�7Ʀ�=����͈��K+�z)/<��0���D�2P��������k�^|y��z���-���р�.�9e��6V��O�&ѳ\ ��ŏ��üoU��G�Gzӏ�2»�ݹ�b���&�\� ���������f#�]��&��{2���1�T��ߋ�W�WG^Lu�-�｛ڲ4�� ���(��͇�;���a��赡��Mo6�bI�����x|ԫ��z_5t̥����Xʖ##Q��z2��r=�t����)i;o�_��,o��
wڏ�|�#1�u����-�sÊ�\l�$�q.pg3Uy����9��<�
���ǸBE�J�!V��.�Cv��/�4�jb�������]d���qy�P�������@$���EI�H;m!�-�ѭ�\T���{�΅Ff�6�tG&�խ>��E�I �(�:4i�嬠2훎+�d�pk��6�U�n�ѽ�Ӻ�dyH�C���0�ϗ)�$��UT�z�_	�7~X�{@$e��̽5YiM�8r�Rd��7H�W�J�g�b�A�/<��`��8����<��]^��"��
!�����)��񎇖ݩ��5R��Ex���ۥ<�nݨ�_��OHX��µkg` ��`�r��/���:�D��p����-:��(�,1�b��Ů�P4	ٝã[�����k�N�_�-�Q�l3�]9�a�n�Ҁ[%�?5U� /`u�=���r�*}���C���
(��x?�a��-Y��>E����C+���&�Vo䕷��T�ya-����8˟�v���rC�����A0~Յ�Y��\u��O�T�sw����l���N�+��$3,P1�3Pl���me��>1/�?��%%]ۧ޲����k�oݑ��RT�}nK� ����"�����lb�vPɨE�v��ܣ�m���S49�7+�V\h�����r$x�P�/ �����}s���.#[r"���gg�˵j'�o�rA��S�zS�g���:c�D�C��2��K���q�r��y���̍f��EB_:��ʶ%�ٗ#)}��|"q�'#'�Z{���G���@�� °<�Dp�
�#ӂ��j"Ӱ�"p�y&E)r�W�%飫�/��Tˮ>�	�&1�vE������=z����KF�M���*�l��邾�%U���K1�	9����1T8F�N��*Y�%[���5$�-,й�x���c�yk)�*Ud(�`dt������*�`!�NcP�?�����Y�ClN1���l^�9'�=G�����66F� �A�5H}zF��e� �
�B�z� _��G�Q�Q~��������G�P�l[O�������(����9�`��,��r���b̓+�Vyaz6��x!a��y����=��ʝ�=E'7G��d?d�&�J��t�K�$� �`ą}a���:��u���������5���4�F�E�<�!K�b��K�B`\<�Ġ�I�k���WPk���eH~c��j��:���=��\��0x.:��iYy�!۩���s3���h�>����A�%נ"�%�����\t|���$�"'�kVY:��I� 5ʼل�T:~��^Q��B�Tf���A�s���qQ�J�%VTb�y�"�ŅI,,�o|7_Վ����\|e���C�T��X�~,� ]K#,	~�\��u�����	�I���Le��P���h�tC�4m��=���vca�ݮ��1vX�� ���,�/"�]������i�iw�}LK1J�CI�>zj���{l������w&�5���q|L/ђ��G��),NFP9�U�i��}HtE�]F��z'��z\��e�nWc����E(�Ό+7f|]0K|tY��[���C\g�Gֻ������o�]y͔X�F0�ʧf����U7V�M�Oɓ���[���	��$����jɵs�	L�S�һ�Og�/+:�0�=��dTʎ�
�/*eV��&��0�\~J
R	�ȉ:TCN_�ѿr��6yu�=�Əm]�c���g��OWL]	��j)`(��[��lI���V��4Wصly�LO6�립��}HivE<����rKjS1���9s�g�Bv��O�j5l�9��69+
�Ӭ�n��q|��n�32� 3�[�XA�ŁKD	D�Q'0�򜩷c�]z}Gde�xO�Z�h�'�٥҈EQq�+�B��Ȑ�Ï�TiR���r�KB5C*���Uzg�<�0Ty5'^��i�:v&tO���V�)���5�pV�b쨗�ۅw�T�^[�ê��qȿ����ڟַ=��k��4��Eg�~��x
���|�!G,E~Y��
�>^P|���2�3G]B (,�-���B���Y�;֢	ke]r��������븞�34�6�^�s�ՃJ�Xi�����n�L��{ �A���b$���uGN��*��ȂN��1�\��h�����2EY\[#��Ś��uʢ���	T�Q�?��#���)�:B�
�Є�� ���p�֢w�@*{���l�; DpH���l���6� j��ofǼ)(���!旧\�/+�S��'xE���D�ˀ��7`�5]e�3��Wx���K$|���t�MP��X��ES����X���i8�+����&
���`�"���Dox,�8+�9V�x� A�ׄI,2��5؉�z#t�4E��*��G����$�YS,�f�K	�q���XcyH���k����!V^H<*�\Ė��G�'k�ȎC�-/?2)�.�51�VR_mqm���Z�$�X:뗓��Qƅo1:2�	���G����q����Hʦg�5�7�h��hU��Z���[$r>���F�K�`�"5�4f��%i�����H���Q"��V{=�mx&����T �b��i���[���m�x��e��T�C�����<���]B��:s;�	�&�͊"�G?Q@c��:�8	k��Zfr���,~�F��<�wG��P��աK��F3�(���Z�={���.uh�ƅI�s��@��fqn�����u�~8�'�|���|�cD<�[/��MN��5��v��s��A.#�F�Hs#������?��3��b���晈&S������?�i�s(V"��h�"�=�������m]�~n�k5���P\���5�Q�^$�,L�����b��3l� Ѻ�N��4�������Ԟ�P��P�kn��b7��axE{�O	�d�>	/��b8-somdHq����+<k��(��^��}�%D��F�Y��Z�?����}�V��+��,q�K���'1��I�%Ⱥ;3oi� ��y�`��.FQŨ��4��]���D�g�~��.$6��wpG���<s����x�˨K����#c� c��EL߸Vd�پ;v1�=|�ۦ���/j*{����M�,5��/�8@�\�t��J��i��s(���ݑ�`����L��*
��%=;˨Pz�/x���^��n���i5*fG����O��hԨ�����cC|���يs��jQ^=�K��N⑱!�s�>��b]7�_S�\�����VS�	�A_.�Ho֓4��l�l^�0%�i�OXs[�Agv��nFp�5��d���e{v��ܝ�$!t]BMKNpY��r�ڨ1�-d�ʐ��_��>'�����0�\�rK%���j������,e������C�_�����U��Z�C�-��k�?Q�_���M��ܜÏ�ފ|2>�B�jsPA�E��rG�~c�,i����~_�Q���������W�1Q�qn]�����Ƌ���$�{�x�����^����c��i�����ن��F�����R�<�@=xg/e�|��6\��̛�HA�_I�#6A�
����Afغ�9M�v	F@q���Cyy�˘>f�	;9�|k
��E�?�hB�ܰ�4AW��*�s�x�B����:�z���/Uk�$���E���H����\���&oM)����|�*��Y��a]7L'����U����Ņ s�-jp�d�ZB͇�|��b������bu R�ku�M�az
B2Wˍ#���	��}+�N�ҥ����c��?8uߤ�o%�d�d��]��{�Qܯ:��h��D�P�� U=e$Y�Io�S:VmF��+�d�:��ȪW��upM^��*Y��-�X�av�E�����۠U;��N*������)��˴�����=���RI�9�&2�`��5)n56��/R�6���f*kH�H3�dD� �����}6�����HN�&g
�������Q��)Y9S��!Z���-Mԇ��8&Ĉ�I��r��/̍��Fy[ޅ�����EK!?��A*����\#F9�C�Zs�b&��+��c�&�#��Y>���c\(`+�`� ��n�=Ԡ(�ը���}��[���T�(��<x�j�s��yc�u"TG2�fs����8Y�l���K)��l�L��!�GSO(*~��W<��U[<�|�7�%�%��w25�Ǡ5��cu��ݜ���m���q��9�8�񆷂ʳ��.�|� �Hs@|��m�� ��dN�^dZQ~�:�?J=�`��!6��v'�{�BV9˅2����I*h/�F�3bؗ��3ӥ�?�@!��8+��Y(�����I��|Լ�N�=�s�nJR=m0��Q"�׆5/�����`�Qh���L;�$v8��wQ����Kߌ��6�jz�}Q*~���}���z�����m�����D������U��1I�ҏ��aw���'ng�]z��8P��`�!�-�2�|�g��Y6'x�Ye��QњvүO���{�$�<cJ��[P��x�w�Mã)���aU?(*�F:�rsG�@8.~��A]=i�x�t��8}���ݭ\�y����3VxR�G��X���� q��e��6��9?����N��f�/�;�J��IS��������ƲG�Lz{K
��`�Lbvw�d�t�N���C����{v�� C�D���p�g���J�9��i��G�#u�����F{ڪb�.l��Sr|�6X	��#͋����ī �/Q�9po��,�Q�č���Ѥ��^������?1.��G(���!�?�rd?�2���m5�4@���L��e9� ���C߈j����2�-���L/$kU�F�4��5c��^@�c��X9�X����m�̧��?�ެ�b��oA�Ne"�Ǿz=`��F����i/? Ԓ;��)@�ʾS�TJ�����%�	���e���/�WE98s�8hS8#̟/a�I��y�x�!l�F�*�9���t��V ))�������t�'Wk`?Qȏs�����z��\g�������s�U�Eߌ>�p>�Dsմހ:��X�?�v����&���ߣ�)�,��o [����f{�g4�)�Tr���������gwD���1�"G�K�*L\���ڊ�d��Q($ꛆ$�oYf��X��i�\6��u�	Ja��^F)oBT�6/kz��Iw�eB�}C7w�h�}ͻ��ٱ�Vuu�ȣ�}C�Fԡ����Q��2���(3��8�4G
rHB��#�ĔXg9p78Xn?�/�<�k6ˍ�K}�6j�����-j�]�As9xdO��a���|so�+t�13�E2��<rȋ�d�Ui޴�E�=�4W��X����?j��Mrb�wAs��#�N��^Q)	�+�׀TX{�y	0�e�<ɔ�E�����9���qY�����XhŖ�w#=>`�JH��TP��;�������"2t���ܸ�-;m
�FT}
xi�A�`�t:.�y�Ը-ݽBk�#�A�sm1G��ؼ$���%�"}v�Z�o�t[�j�«�ʡ" ��jO�b
|�y�)���߶�l���+���#&�(��b���㴪�g�s�%ɓ�����d�]B@֠ z�}��ۄ�!��T����i��"ȉ=K c'�!�(��>���}F�AXDь}�4��P�ꌓ�M*ɝ���X��47)3߲��2���IfR��?DH�&IM ~�b����S_n�F���m���*��Pw��(�k����H������R�.�UApLo�f�i3A������{v�~�G�DV�<�Jө�ż`�Q�t!��+��f�������7��X%3�Щ���A!��X#��E��h��[��5%5$��#9ؤ���j�xbR�����q��n�ܬ��n�VR��F:�
���J�W���\�Ϗ ��^���B��V�Y2��ǳ�����L��'�/ܘ�6f�Y���8_�ӛ?|Ѳ�C����|�YbE�� T�%WM�J�<Bȭ��y��#��?���(��\�����@lX�`���/'>�6h:Se	�a�/�߷�N�.�|~Qy��H}�1#-�Ʉ������L���I{�e킶a�hq��ٜ9�H&��-�����s��6}F6x|�(
�P������Y�n��f�x�˼U��7Ys9L�.P�w�Z�{:ѓ�뺄%i��l�Ё@�(�ݘ p!@��ke�qg@�P�%�K\����q�ܣö���D&�ZRU��~<�t�,�c��G��ѷ*���V�y�AoU
j�-[������qS�3�\�v�Qhr1�!��&l�G�����,���ܭ�s��- �
�8bm����z���Q���y@cU�<]έ�Wpr�Re���#.���>q�haL���
�����q���Ơ[�2��B��k��@fġ��f�����4jZK_*l��(E���3����[U�n	�q��(�,�`fLu��IX�ǽipN�oH�^u������Ag�����[S�q>�Ӌ<���?w�-@�ZF���QMat%�������$s8o.�ӊ�y�;B��'{~B��_��a�7Ą8��h��`��I������Bv*�	�C�����@k*�����-�v��?�S�'�r("p�/��v�R[+U+#�:1�l]�z�5�sD�9'E���mA�@��_~Yf� Q��J[8h�	�&癟��'�C��d�2<�)ȁ|lk}�w:<a�I���G����˺��/�
�ǫY.�����\n��7e�^�E4r�T�u��0"�w�l�_
AJAS�&�5��U�&���U.U��+o���션��>��*nd1���^|�U�F������ms,��GPa:��5���[�ΰ+ջ]�s�eG�:�Yq�$� �EY��"�t!	:�(�w烓oln�3	���}�IXˊ�ǭH�1�K�͏�q�=*4b������?�����W�C�	+�+�,kl1V�?���:�S>[�ؓċ�瑈�.��bc�s�<���<=�yΜ��O�OA�S�[����(\��/��>�	�
�l�&PׄIS�̃ܞ��#7ʀ�{s��X~����%xR�jF��"�`�ek�U_�9�*�1��5sę����l^�zO߯!_L�d_�@D�v�oN�*$7�lŞ����w�	��a�;Y��f�Q�L����,�����4����K���Ҟ�����6*ٝZ"ը��03�
��眵�63�4��}����/��$��}��3����h��|=����ԩCF�B�-@�+��a�Q�K����o�`����=2�����5՚���S�O�� ������o[@[0�*�g�\�vx�L��4j9V��袓��N��"�?7�OOH�A�ӑ�߅*f��bM��EQ�qΫ���(<���(��!3|��E�"e�J:���?)����0q`QY9n��Ro
P���"Ќ�ɘ��|!=�����0ab����0Z��wZ�=|z��w���w���`�}	����U]޽ܥ��2�O�2YCb��g
��%e#��Nû�|�>�v����\��R� �9?�
�B��
IE���V�E^�����bU���s�cd�p�Z��{fj�G�P=5n��%zŉ��cG8 �@e9��/����M@��SPC��'�8]f�y���T/�4,�X���|ٗ�f������E�6�z�0��͙L��ꥳn)��~Zy���WM����qHoua���^J�p�ޠ�~��1�s�����x<�=����	T�08�ŀ�A2��e %�ߪV��\C,�.�Ȭ�PV��־(��f�.;�.S��¤��da�\J�?L'��LvŅ�Ɏ�Ӵ��,�i�N�e\����Z?[�$8�R��L�q���ʢLC��G����u,M��%��0&��mȓk��M	����|�*q�D����D�lw��fce q�����э	`�[j�2*\��@�Q��<�-���N��� |��(�Xf���/����q��>w�����;��v�"���m�M�-
c}�Eg��:�`Z!�`h8Rv>���@o�H����]?��¹�O/��W�J��E^nc�&X�ڢ�eV�U�~x7� ��r�gC6�;<OYQ
�W_�ڻW�ʴ�������]���D��R��.j��9<���I����I�D{���+�]�-���<�	%B�6s���5�0�J
��k�u.��9�n֞�����_�5OOn,D�벧H�䃶e{����e�"��H|�/��q�6������ݴ������;���*��2Y�~��U?%�A`�%k�Qb�Z\hlI��1��_�6鞑��3����R���A��ږ�~m3D�g�n�#�v�Ǉ��(���o���1wv~�P5�ؐ��Aڷ{"���Z@=�Y�P�ԍ�L	�_ٸ��0��AWd"���[�U��	�W� ���^�3j���hń֖��Y�a+ό�Bs?��p�lWG��< ����J�7��:%���Th���`Xy#��W��ȏ�v5AXJ�
ޠ��M�Ӣ����)�?+E����$��?䟝�*�1u�B�-��4Na��!�|�0���3��?m����Zג^�]y�z��XO�swZ�b��K­�!�nho�:���^:�t�{�J�D�xGEպl�?�v�3���e��d��5yA��A�����?A(�r:�bmXT�}�Y�6��Kή'��k�'\�%ԘR��F�?A�n�X��V����U�ه�֮:�S�l��^��vL.-��jS���9>0�����:������#�D�c�������F.��A���T��yi(T�L��H��R5�A?�EYu���P���q�#��0��G��Jd����;JS~�AvM��<��$-H�� ���N�Ƕ��3��0��@���	"f�ƫ���qr�G"�%���s���͉�YLն�&�um�����,{�3f �:c�?�n�p��d���j6�&V���2�����D��d��dM���ʠ]���1K�����?����{;آ ҥ�{|S@�y�I:댱����6�Q�L�2]���	��,�Y,g��$�i&Z$}�R��k��z�Gz��-"��ÛJfS�%f#}@$�U��5�	�����o�v{��j����DX�shμ��ںhc)��*o��B���l��e�U���������8~?�I��8��g�F��J�%~��yP,\+��^ٕ��M���.VL�Z�V,�y���&�h�۔tћ���`�IQD'<�_&���oY��[���Z��J��=���6B7���M�,_�6�E�^�r���Gϔ(Δu���+k# =�㧭=�g�`�/1��ô>u��Mn:�h�'S�ƣ�xiWY�b7K��B<A#m���};�a�
�Ag�~Ոi�႐���v���&T��3J�Pp�C{���	���<����.L2$����0$҃��]����-5�����?x�ī���jM��������M�Gw�~�S���Kye��S� ���x�\��:����N���U�����=����C������ ����q�b%�\���3�^.��� {d0+ȵDF4r(a�rU̱[�}�p��C�8�m�eޡ(F����7�{2�W��b<�r:�`�Q�@SƛyM&�׏�K���GUλș�	��Jm�AP&t�&�v����GQ�rS���≡������ipҸ= ��\7�>< 6�8�zک�,_��8$yp11��I )�B�D�l��^=����*X�$C���=V�)��<���L���.��epzQ�ıL�9�g����&�e���-a"�R'źw�޷�̿��t�mQ�οK�Zo?�������*��g2~4��t�$�h錦��
]����0�������&���`��	��{�z�1�!d@8(�^Y��H�:�5��8�%c���l�@�\o�U(�-�^��{C����t����&ЅA2X?P-�0��(��/"��}S}f7��x�v��9~�����SNA�ջe:�T4	��R��eh~82$�Ǩ�VM=g",��LW`ݐU�w7��us&||�+��(u:#���f&��z���K��&8�rjRm}(���b���B&I�������t�����#�؁�$4U��� �M��S���g���E��%�̒���3I��T���{��-6fS�!6�ť��9�
R�`��!f�iI���-~0�.^�	���!���?��/k:����"���W!��g3Z�҇��b�@YV�\h�:[�ʧ�(qA,�hf�e��\	̛��m �G��3�S���{�+K_�b�a����ֿ��	m�ب�|LBX��_��)��j�:%!��Q+��\+<ݵ{�����B�Z�HK���v �r_GV�����0x�g�0���:��keT��*�,��A��B��1+N�xZ��Q&T�v���H&積��Gu�R��H�9W&����g' 
���Kh��xa�w�:Sǥ7�E)�B���r�ex���9�'�i/��U6���d�wu�\�"��	-���y�/��RF^!����C�q��[0X�\1 '[�*�`�CsAдv�quE�N{�'j���a.쥿�㍛�����)Iҍf���~^Ss���6]@&Ǖ;���%1�J���V�w��C �}���Uף�t���5��,��ҸQ��Be�驦�Wm����"��!\��z��H��h���r��>�����k��Dx�>O���	�T/�B���eG(�Е���Q�Q�הxʻ	;�2�z��Q�*~��WN�5-��zs���ϥw˭�:�y�5�>1���VJ9lo��GĂ[Z�ˍ$�#�;`��2H�$Z�&&l2�!w
���l���ۡb�� �|µ�����c�~	ZJ��a�+�.�[��q'�����D����,	��`X�E ?�`"n�ӳ�P��zN �k�T�s/66B9Fʊ��Ν���b�|&�I�^�	G猃��,��U���80�=�$��6�(~L��GO��Ѧ���I���J� ]y<b��DK��kO,����!���f��\X�߷��U���A%�g��g$@�D{�!��_�1�"kc�]����ϲU�܊O譮a2[J6o�^T����ܒ�!]��ݒ���o���Q�*��������u��4/I�n:Sj�M�c�>���d��Ϻ�nNڸ���U����p p��'���|l��_�^�,b%jHs�iz ��ko�:���SҤ3��l�f�ӭS"�!)V�D7P�9ܸ�b.��Ч1�`�5����I-\�{튱ڨ&�?U�����NO4�~wM�(vd\�V�;�գ�a�5h2�%X!�W\���Ϲ޿���YF�������s����	�S)�V�@�j�i�CX��E�紩Ԭʀ^����_1�㴽ӈ�*�����c. �6X/�����K��+#Mz�1��"��(��P���9]K�_��������P]��)�}�+�Q�?��/M�	<c��O���{��`��7�7|䈠	�}y�?���6m�3�����
�x��Z|:��o�M>� �@�#/&�����/�q��@���}��_I
��{>�ߪ׌N��r�q6�����j���"�3�� j�}�,s2�װ�����ۻL��C_�d:�K\� ���@}�jH�`?�5��1�FI�@�Y�A�� ����sM����P �m[��M��7�|�{��@4��c�+`�i\�0OD�ς_
X��u���jYR�U.�z4�/�3&>�<d\ύv����d���+��È�"������hC䮢��T�raT�V˺�Cs����Gr��Զ�,�5�t�>�A�pÅP]	�����8¼=9���_�c���~6A9�Q����!�8�!�WC���2���dp�"�s�|T��93�B�O����>S�|m� ���ޚ��ٓ�bH��rf�����"n�)$U�P2��|{,��F���x�!�a���;5�g�8a*�:��5{�Μ��x���_�-�B2���D����]\�z�s�`��R~,�[�D-`,���u�����H IOↆ �AҤ��33�f���J�2x߻4�vi��j��̋����?�rݾ�1vG�J�%d���!����q2����?�|�q�2���0�n�}>>a>S�M`��S}�x���<�&Ќ�MO!��"ت�	
�����<dE��f�^��$���do�?;�U���i�1�TŰz��ӊ9���Rl�^�E�b�F�����m�������TL��\���ZR���?e��E7�ɀ���:�V�j�&#q��Y��� E��+CU��7��6����Cǀ`u~� �7�y�$�\�zŰs�2ѝ��.�jg��ۨn���,�|]:�Q'ȯi����F�@����\���ӸFK��Q��%���u����O�|nJ���0�p��_�����M-^����C��~�(vf�R	��(�r@i�Z�l�URcF�@�/@Ua�!�^��cD��#�c:��e�wٟ��4eq�E]h�'��Q_l�l��S��ŕ��"[X����ھ���ò���~�f�6����?�A���z�(6M�ĳ2f|~_�0�0Bx���s�a'Ӿ�N�s�^��ܿgd���i���%��Z,���!���ž���n�G�0B�m�}�_F�s�L�5lR�I	�!(�M;2�,�`����ZY�N�d����]�'��G��Q��s��F{���3��I0������ص��q��5�~B=�C��~`Y�\�e�Df|��˽;<k�5��=���/u �rju��as��2�Jd7C�T�đ�|��a�!X�E�ňNtQ
�_����Tm�^p��"jdg;$V����q`y�<���7|��"��?E���$.	J!�g"�?��(J�J�����iu�D[��ഉȮ~C�I�������ǆ�=q��.dU)iyVNt+�x�B�˨��[p	�}2d�%-�K�#b�G)}5�UVX�8��V��h����2,Ei-�~BTc�������8w�n�S���F���4�Y�����o�y\�S�%�IpO�T2�0.�綶{!�J~��3�|$�Ύ���30��p��n^-9_�p�/ȺXԛ�v��)�
w������[�H~x��U���o�m�5��B�Y�U)�|�p�]^�^�V���y��*��f�D�bJ����J�,И����O=����*�����'8��!M8}���V�@b�3�e�E�HC��yKƲ!(2R]������jI�'��EE|y�1�)�3z�R��O�2�0m`(�ŖY�.��S桠�f,Sz�Z�o��Z��5uO�8c�kk�_���ȇ��r�6�n\�@� 7���a%f&������L��4u��Ϩ�Wh�J��9	W���=D�����*1����� �R�=�{����</���p?}���$��f���K��D󓰱`Av���V�v���3�͋�7l�@%�'�����e���+�!|i��T��r��4:$2֝Uk��l��σ���엖���kmN�W�`d��/g�;8t6�B5�Cy||�@>�J�q����l#i��'��	p�F������W��giT��&ٗ�/|���`<���� ��މ�vD�4;��{���x0�n���{�Nu�ܢ�1�?b�����h�R§�M�p��Ls��)C�@���aa��E����w���d����Q5�f0����k�zø,�����dO+=�xDd��G��&�'��&�穔"�|���;����r���c�;(��BE�r>���QJS����頩�ra��WN˵E���`��ĝ���"�ʁ�j
���L��<җ�36�7}?l�&
���\�3()��l��N%k\ӟ`���|2N�~�\y�����Q��0F3���+�����/��K���^��}V�R�q6�ͨ�V��K����Z\% {�͆�.Ϧ�G���LG+�g�Em�d�U������#<��V,�V��[�Xe��v�@���!�P��lVp��:�.k��ҮP38~����1#C�Q�\W8���1��Z�[��U� ��6Bs.�û]��:lði���_� �1��D�,�i�o�"����M���3�}:�E��Cq��9��c���'�������B�6NL��Vƫ;��_؞� l��,���Ժ��\^UIWH��Ur���6��]�F������l��+x*�2M�|��68pe��]���p�!�St�.����V��#x>�2*��R�{�߇u`���,��'�P��ľ���(�	�'�	�44������o��Z$�����%��w�1���IqufKp��XV#���,{��Bſ��J�~}�S@�'��`�m���:Yy#�LG�W�`/���4�Z+��du䈏�(㭪�=q�N��	���Ft�ش��~ƒ�P�e�w��I�q�٘����EvN��Y��g�rq��S�ߥ.�S|4�86���i�t�$WC^��NP�a�2��F?�fEo�P�y�HT���o�I9Ҫ��s���'�HX"f2Ĺ�[u%5�|Y�����~ke��Bn���a*nӃ5!Ey�``t �U|�@?Lε͚��8���ң�r�v�o���>�xxuZ�o����r"���C��ތ���ner���U�B�^.V��<�fFi�P��蕯�����,��8��s���{jv��@V!���i|0n�@D=��7h�t��,;|R��Oרp_���7z"�V�?�Q��4�/�ɏ�=ߣ\����|a<���n}׸�?�͌O=�R��VM���S�V̉�Ӈ�F�Ʉ��N�Q������* �*�'�s�K>��ϻ: �|(��Oo2�`0�RA���`�TUjee\��>�߲����B�p_�Hy��
*n�����Π���� �f�Mr��x\؎�l�ȼK���O�;Ӊ,���������s��ŋ���Etu�<�4R���7�V_��J���8�*��	����\���b�p���Łh���,�9+8���{9
ZK�c\��`�oZ�b"W�?t~Aר�#�g4�A���ڈJ�+���M��%��S��Tߍ���{$�]�$�qYXЈ���MS�sT�&ZX�]��n
ܰq�0�ԡ(&'PbC���v���O�Y����j�_@��藓�++sU	}h2���z]���|V��NSRG��^>�8�{x�E�|E�H��>�ӆ\�j����Ů��#�����vzb�'�l*��	o'e#�*p%�^�]� Q����>mR�) �}��A,��)�h���3�<��!;flZ��� ��� ������S&ν���:rYG�ӛC0;�����3q�'�ڎY��%i�_пXe U�c3�,t֏M���Zv�cK�ǅ�/.�1� �[�����(1�2�3�Es�s�	�烳��3E²�˓�C ��X�·�b��]����>.i6��"u��b5� \���֕gs�����$L�w�k@�]���G�d��Q	�3I �pu{#�D}�	m�J�x�Sm�(��������W��pZ���&�������H�W�g�ı�<a
�:Jv~O� �=��S��ק�2U-���S�[ɇ�T�D��耡�Ph�=↖0�AB�yg�"|9U�w�6q"�$xͷ��GHk�XO��� \uH��1Im�U�C�Db�Խw��{��@0c �q�EA
T"��V�5��1�>�	��g��iPl�e @%��1$�v�`�P�u�X���;��L�:W=�^� �m�V`��	Zx� dLTγiϽS|�)s�u}��0j�ak#��x��_��9�fC2��u&�:(� ��t�t@1^Ե�5�[9�u� �7(���G�e��?gkl&����)(��7���tg�jt�T}xn�4!�&\��-�i����~T�\jI��
�ж~o��KTl\�����d~~e�-�>t�WQ�{=�T�Hyc�,�g�t�7(
�1�*m�ǂ��P)�A����u����Z����Z���mݼ�%�uF%~�9��Z����t7�Q��
�4B�ZD�%z�;L�e�nX#w�zS6�ln�|�Y0�>�5��V��BȑU�*�G@�1w��g�����f�4���emx��٬/y�f;� �Hty�]N�_���"_��?wC�� x����i�v|L���m4U��7zE�V}Oq�P�d����8��.|�9�����?�F�������k���VQ}�w�ow*�Z+uEڤ|�@ �Iu�H��U���{#��L���m4��4��M
B^jGH(ǚd����4�	��>_�Z6vK(��tnOfj�^��z�>`	�L0V��2���*��׫��@�T��S�2��j�qx��P@�����y�RD*E��
�1{��R�)i_4_����E��ԒY����Ӛ
���k���i�b9�T�����d,�{��e�A���eq�p@����wǄ	G(��y���Kiv����5����Y}}:y�E�ڢ)�V	ߧnD����/n���&���V,R��l�P�G��HH���
k���Dū-�o��i�|��jD���"-���:rot�}�7Pc������X��9�$�W��V��X�n��Mϗupw������B��.��lK�Ե�fn�}j�$hx�h��1����k�9N\���f*�`����\���{`��j�ײo~>'�T%����~�����&��Hڵ�\��n�1���NxX�'ߪ/c��������������p|���&�Εa|nS��2buʭ*��O\2����W:����S�K
��������AA`I�l{0���d]��jgj�V��^|� �Q
4W��^{��g���c,%��sQ�x�W߆��>��-	��᫔S�_���7�Ot�|��ɉ��� ۿ��@���=e���,��'�GF�����XǸH�'3P��o��/S����]Y#�)�ne��:-�8���ޟ�ޭ���U���*o�C�])T�d^��[�BK58ˇ�hf�c����u�-�22��v�q�	�A�3q�3h��T��wq:���Ԧs,� 3����d��� N)���i ��Ҙ$R�?�:��7u�jXg�(��� 9��K��l���/)��Ñ�_�@��?z��M���k-��c+m��J{��~�$\Iؿ��_��6��I������3��Z�~���d%��F��5���;����V+��M�7Ju@?=`V�!jf=W�z�^�cs)}v2~���:����3��,�yP'�>���y�b��/kE�ۂɵ�^���VH�E ���֪;l.��2�q|}Ko�/��F��u�F\��<�7���X��sƱ��h0����(#xH�Q�i9�0�6M2�;q�5�j��9�Rg�YJr	�b8��v���b`��)��51Z����Ĥ��� c ߽E��	�;e-iO߉�Ƕ��7T) *�x��I|7�BNu�s�W�X"9�����Jf������%��F롥S��E}~�C)�L)���m�}���4L�K��kH쒛($����Ň��r4'�,y�§0ͻIޑ_�D}���85�L�������e�L�[L+�J�-&\�{������Ӊv��Wlb[���̤��u0N?��	����$�fj�~G��퓵�C�����Ԇ������(+̸Lف;Z}b�?��_d�e�z�Ԝ3���%acy�(u��^e(��aZlc�f9=��C2ԟJ�b�ח3�ߎZA�^�7���J�����-��~Z!oR�@ʶq���"6��R�崕�C��uJ���W	���͝�A���G^�U̦d `�R)�e��A*X������8:��y0�|~���#{@((�p$�xsHGKr���L����_
X-�����d�����l,�����V������D����
�ee���¾�P�?���agO>_�wn|]q��Q�sYέlBDK$�@� �Ѱ��A����y���I��]v�+�h�$���oʒ��>u�rx#@�Q!��Ѣ*	�Vw�E"�ʕEK[Gb�n�ھ�Z-ǟ"j�g�u1	y����w6U?�&���wL�ۯ�)��Y/���e��
}{�2��Pb�B�">䠃��18+��:�Tr�����6m�!e(% f��K��$��t�����\��--�	�L�ˉ��W���@w�Gj}^�V=��U�k���ԣB�j6�v/U	(���K9n�=].xI���5���=�t�}t��(�p9�B^��D|J�10�[�74ŧ�i�?��@U�?r�q6��cR��&����c��V��0��ɏ��a�stL�%����"J%�����Dѻ6C�e�� u����v�a��;��q#@s
�X��࿹p���rRH�T���N&����� �v'�-wyh��n�-�{<��}M����h��DF���h� �i�@#H�� �a0ݸ}��M�뼽���?sקT���-:�Vw{���8��,���ڄ���#U�0�8r�S�%��yg�lݗ0g��(.͍��в����N�`�6��P��t@�#"Xn�A����:OOJ��M�@5���Y�X�2��-vc�o6�U��9�7���5�*���Vͅ�����7=oy�6y+�����f�g����ܛwl��/��4*N=e�Q�#sǥVX�G��UL�ٵ
@�9z�31д���Ņ�wW��X�~��������2A���XK)���ų��w�sX2�g�]<f�����C���Gd�6��@�� a�u�k���n<wf��� <@��S��rҪҰ�x�%ved@��B�%��X�����e�;�(��͖��3	K���@o�:�Ҏ!� A
�C�N�ְ/���S�Fb�p9��k�LI�z�uɖOa���{���B�Y�gE�Bdf�ؚg��ҁe,���F��v�C��F�P1dDP�}	Va��]��׸u�h�į� �^u����@�)w��O��⤓Q�$�88
���էY����4�w�6����5iL�X��E��7�|fu�3�d�O��ӷ6?��
���}+	�!���N�1�4�@Mgz���El��1�
PHSǴ�<k�T&f��f�r���D��)���zgHF)���;ń]�&k�Z���BŁ��U��+�Ii�K��!�}M�P�0��vN���>�LhknJ��غ��C]�/=U\bt�w�����ll9[*_����KKy&,dڋ��_�q�R�~=���,+Z@�.�E��-���砨��Ǆ�?���� R?�,�*�z������X+�N",}���/��!�P�7�~�ӥ�,X�b~�|Z!wdW@�K��
,��֜���p���H����U���|�<����[2r�.������<j�Q
�or��x>�j��K��R��"�^�&H��M̭�o>�������7�53�Z�鏑�]M1'�̍���0�w�[8|��6��7K�r�����C~��TCq6����C`>�%�0��o�����[D^ʐK��\�T�C; ��Cu��-�bO;��$/��5�<=o.%v���́�*q����	�2��:�	{�l�p����д@W��k������4&�S:Dhp8�[9Y�%[N�|Oً����OpB��p|�&e�H"�d'z����p+I�������ZP��+�]:�\����X%���K�'��L*����Zj�+=7R�F�,Z�"�?7��\p��3l�r��\�7�������Q���~I�� ��0�o�92�!�"�.�����}~->�l��T�&��(4�a�o�q�";"�����%�]Pj�"���J��bV�hu`��]Y6R+����J���|�'���ZBe]�-Z��9)��������գkQ����ĺ�.#Y��f�:�;�`�āB20&�Q���!,��Q���dD_�� ���S@����rk�T4���u9t�N��EmGH�x��o��63�w�;���)�L\iA!*b^��K�imC�X1֍�]�2IQ&�c�'�(��?�0A����Y�"^9Jе�	 v�'����>W���rb:�p��ĳ��		X���M��+xH�ɒ١V-|��J�Z���ޥh���)v��yg�}�&�+�RG����K+���M�FcH�%W�h���e�����8?��kU	IUR,/��[�A>a����ZOY��Qp�G���<��֏a�k�5��?k ��>�£<oZ����"��r��S,�g/r6�~�Eü�=7��E���;I� }g��ԇ�O[�-R��`��#�
d!1[�X��"���]�2!C0O8�4�̟.�Ao"p����}[�����e�u��j���u�Ӵx���\�]0�&�����\^��=FPvx�M&p�xqz������n�^9�KM�-h�	��2Wτ$��������g1������ߖ�|�Ft��ѱY�녪`�S�9�\n�?���r��*>���`H��E�;�fP*\�8!�U$�Ɔek�c���j�iL�[bG�.���!_}x�6�[�&�e�{0㓍����cF��qB%yL���|���DN�R���=ԉ�����)�[C���3��� �?T��:��ө�9�f�G����g�\vHQ��SR�9�4�QLi��۔�1TtRys���eRSGXA7�ރ��M旛�<������$[=��q�J��B� W��®�Xm�т��\�y�G����p�{��My���2��sjD5\0o�-.Ɓ�G���D�g؛���F^+W�t<tx+����/×RlS;y�,�Ϛ��BgQ����C�H80)�=&U��\!q����,�p;PR���)cI���y�C>*X&j��<��J�
H��`���N�A�yU7�9�
�<2�֞;��o���1U�fYJ�J��rӪ��,j��),߸_ē����;˻��i�Z�YȨ������ܑQ��=+���9��	:ORm��Χ���V�[	t��n����B��"D��\��e3ۂ���!��)��h��v��nx�ޱy&H����S��|&g�j��$��tǥ�<���e-���z�i�T��Gu�H�����-g��[J>r(�0b�*ORCm�ɫ{�C�0lKRřh��?3�F���Ү�[��=ӱ3h�8��������+�H-X���1}b�'F�#-�#V7�:��rUΪ9��B?|#O_�K_~��CcbS�[��J/G���OO�8��]=�
5/+:�@0�G\b5��/mɵ�+���	�#�}b��uV}F�v<��h�!+�B��E(����e��	�>�C-�g��I��t���qB]�Ȥ��L�$H�ܷa����0 �[���$����+�����$�t�,��ʼ�">�Ђ��L�b0sY�cһ#��<�-bh�fv�]���q�i�p/vVߘ�m��r�A�\��#�q�	��(z��B�nQu�ذ�e`&�M�RI��Ϳ���s��?�i$���Q���} T��b���rn����i��.'nB 
 �۪ �j\� ����s���h ̚������4�UC!\�����t�׍����=�>Ϧ�di�o��G������q>�^ᮃy$C��|�)n�]�A]��_��h;�F�9�+�5VB}���,� gًR�� W�4�բN��1�$���
��	TJ��8���Q�� �G`d���1��=!��,HN�^��y	{�)�w�ݙz,�`CFx�3�J�kFL583����H5��h[��\��"x)l^o���P��rp4)w�s�tNEu�y���mhc�L����F2k���@�8�V�f�S�d�{2#�<	���~�� ��Q��ј���<<�Z�O��>�8ڿ�b\����(n`���K�ɻnx�l #�y������k��QN���o݈ؒ�����<�����ӷ^)<=B����w��)9	�dJjl�E�ZeG�K'���<J��^.P�%�̖u��AYk�����/�c$!�a҄!M�{��K�A�$X�JԜ���~�������m��G��-�q1��g�e���>3"$7�`�L[+?z�c�`X�݌
�����\P��Gy�qf��ݤ'�ru	Kwy ��I�,S��-�\�.���~q̦��Td�x����~��s�]�F=|)�`�P�f~��M��)2&�o�e�L$��C�č��˺jp�6�l�%�� }ƌ�a�5m4�6����%߈Y5,��?��$����\���7��`Nq�Q�g�*l9C=�f<��P�\�`��mϫ�F�85����� ��[���q���P�b�ӄ}Rd0�i�l���r׼y�ʮ�9z��G^A���<�f��8������*K*}����!���W�3�D=�6B�Žp��*���^�f�ڿ��[.CQ����/�d�U�bŉh("��d̀1���������ȾzͰt���!��I�A���>�2E�Ǫ�۱9Fꔬ�W��fk�^ףN��?������(9��tZe��7��"'5h�w[�S�E���Li��ݓ����;��c�􄅟0¤�N]�$t��	&�Do��ZK����݂�ᤧG�)�N^�	��%Jd+0)�Eƅ~�W�"O�m����F)��ܼ�jO`��G���^�|���� 5�cS�Ij�0�SX���J�Ñ�������������Ih!�y�.� ���o��JB�f�J*�ތ���+� qf�
W���U���B�����я�����k�=�׊J�m%�	f~ߤ��(�HJ�0��v`��饙�d��P������F	�ח��2�vt%E�F�4�S��o��N�V���O�r����)� ��������Fy��՝�<�&�-uh�N�ol��Y2!Z���ǂL��#�9ʊ��1�ٓ��jF>�j ��b�l}/�i'��p1��A!���j��ڠ��/��z��b����	�����(��z�x^�������R^XJ~m���hi���:�1}�=ƮN�$�n&����⮙<2�-�>�r�䲮����X��Lm��	l��K��皅�(�-�ȣ����I�"T
�}�!d�$��N�q���/��I=�3I/%mwD={[����� k�CW������0�����<DɉzO`PT��4��0�I�����=\n,�K��a'6����wu�ہih���.��Ƿ�&�g>ȸ��l���h��Q����|�EߞZ�:��{|Y��ʵ��_�H�0�ks"O��| ��D�G#29�qڨY�^���̎+8��y��R������W�*� !پR�����
�T`s�C�2�p^���79)�e�oX+����������MUH�c���I\!���A�5yn���#P��j���iWkT?V<h%��Ppw�"�6��Ĕ�u��)�KM��������횤`ɺ ��22�Nn;�j�fSv�e^M�oc����*�3&g�ɜ�V�&�=����v�_*�c�~u����L"��v�23�\&�C��\y��e��|��F{�W�~ԯ��-o��	�����ohO�j�&��6���囈������ՙk��ⵕj4�m!MfǧKr��G��i?3,�aG-�W������Z����ʶ�1�+-�[|g�� ���Kq����`�J���t5��>��Xމ/���, �fd��u�5�n.Y=�+����4�cRt-��{��#��䲌���n�^]�6�Ia@K|*�ƺU�k��Ly�3zJ�#zR�Q���w"0-�� F������!�Z����ư�n�����X߇��ߘ��R�g�}*�}Rᐴ��q̼�R�?P���ΜQ��mW�/�D!��žr'���]�v�kp2C�d[����;�4�S���{/~X�o8J�U�.ڔmv�7��� ~0L�6%����`�F�h�@.�[��)9x^�������?
EoE
��W�qԇ�tϒ.Sd�S��˦k��L $N� w6Rx��~j����S�>�~&��K�޺��]�ڟ�t�fw�@߱�4�+8F������!��Ȱ�����>H��\ N �x����HT��uq�ҕ/�/����x�xe��ojk<�btɃ���e�~��'����<:��N���an�-���A����x<!��3�
�@[P��(��E�y�V�2�$�j������&��*�HI_93~��_��C݄���@�o��I��S���H�����>.�v�S��������<�PI��n�'lVr{P�~<���gj�o��v�V%��K���Eq�m(�F8 U�N��0;�+9k�%��w!o�v���5ʋ��7��K=���|�y�(l��D҈kBy����p�uj�;q����(���`�А� �Ş�����1�Ms�4)�Y�o`g���s��Q����*y��D�;-S��!ҳN��w��{IU�;{��Ũ�Q�J�ZI�N��=t�����C�M����vI�Ƶ\420 �+Ѿ��������t�-�TKVxWS�3�]���~���T4E�R�b%_m�n�]d ��h��KA��q�XK�c���z3{��s�>�c̑�hy����7�e@�$i�`�G`�:P�����c�:6oi�����@DF��@{B{�lαC������8��thžirIx�"��&��d{�K�:���c���W��!?l-�U�'��?Z{����F]�Z{�}#�r�R�K�G2U�uIa67rԋ���!�zU�(���Fw<�'T�\�1���Sa{\d�4)Ў�(�`��tL��	@5������d�/�&�x�����}����`lB�W?��իF��WLbM��X�/H̡�4���h�0�|9�;����gt�[T��w?x%H_������������p]�1�jQLI����i���a���n���*����FS(�K�v3N�s��@�䇓�|ˁ��"����9����uiE("�|Q�$MB>�+Rv�86��b�����0�B�j�Q����NH�]Fw���oF�0��aT0��r�6��.U��>�q�*��Kc��e�/]�=Ȩ'�wM����@�Ex[k	�o�h8�E��#l���+�k�}$% Z�rZ� �m�8�x9ZWv�;�e���������y��X����Ct
��\�u�Y
�}J8�|�}�ܖw�yZ�x��Z1Zw���]���P�#���i��'�)0�>��t�����.�����|^*��/�luׄA.8}�*�.��:�e�̋���\_eN���э�߽��G�&��48u��FEj�����R��9pٸh��
|*�f�^�\�8�y��q�.�3R,:$��x��Y�˩N���H��C�y���Q[KC$��&�t'Ԓ�(��Ea{� �[W���8&zX&�����^;��1}��~{��'������I��u4��DZ�Sm�Q�FY���j
)hB-��E�)Yw+hq�JU4H���.��iu�w���'جĆ.�(6@X�!�X���GJ?5�Ɵ����>נ?��Xkx������̑Ph!�g �+1�>����~	R|�"�Y\���~個	O�C��9P-�	�c�q5X=
S
3��3�����c��+S��]�I����\�
�\Z���T����B��A�qغ�U�3mj|^W�gyׂj�9�;Kn����{i�m�?A	����ys�`θ�r�r���FۓKQ��d�6���L��p
s�S�x8��{�\7wkn���.~���3X���v_�p� ��(�ѓ�*�T�1�l�taN��@����b�*�ZrxAj�P�<�r>r����b�gk��1�'��4�hv���u��־2��

l�≸: ��R:ʋ�A���;BHr,���-PRk)�ɘT�GZ$�&�:�U�zU��a� �N2�1A�����3���A���8OP_Hi�y "���o5L���aN&!�w�jr���i�C�ѓ�F���$\xf�Crl�Z����S�}ïnA��B�v���_`���T�`���~v�w@j폎�Y�j�/r>'1�4]d*��I-�j�������}G���E���3��G���s��0���v��:En<��wt��l@�)��6vJ�V�k�Q�p`�HiBX����v��C!�q�iHd�������<.k�~�,&����R� �b��� ���>dY�CY1\�4�cܴ�̡�O�z�S�����/Z�%�\����y�&2*���Sm��҇�}��2���q=��N
�ݨ��r��9I��M�����&���g�e�k���^�{k&�7ĕ5�Vd�I��L?�|�K��݉(���^����ib�̟��	^mW��Z�z�AX��y0�ZI�{jK}/ъ>T��h�6��	"L��k�A��{��25�����!_p�}؜��b���?M|W�*[�ʨ(��# =�[5u��=͌,f���ug3�蘖����.�Jn(^��.���C���py���2���0oh��Ѓt�M�4:b.1�Cd�� "xb>б�.dG�?�=��S�슻W��*��
�ť`���a����e�������c�_�"��O|ϕ�6�u�&܊K�vi��-$�����ˤ�ay�HQ�r��� ���]�5���&�7D�^#������s�i�2M�ǾC�ٛ�#�l:��6>����oq�S�W�+�Vk�/�A�&�c�����{/��� ]ov�w(C�WH�� �6��a��x�w3�N� 4���W�'R0�÷�E��恩�Jj}�N%�����Es�m��vEZY�%u�/U��k��_-�������FT���f1��T�s��>��̩�2el�!�FΓ�3���`b��W`�hɊ.3��Jн��r�D~��[-'�֫zu�#Q�0��u[ـ�UG�P���p�p)rʁ��*���*M�SH<@i"��`����r�z����?� �0�9�9��LFr���Z �I��n�,�R(f͹{�����;n�VWpF�����/.d���%,;���J#��+=F�[p��Pa-ZA��Z�ۀB��9�o�� 3�J�WAX����>a_�N��kL�}=��/>ds� n���8�慌��D\n-���>ܪ�~��95���y�U��Ec��Y�b᥄�`*���'���:rTm/�j	,��x�~�=]N'9��Yԑ �-1�W��;�"@<�@��,f�Ш.���}{�q+� 
�1�����`������	�ӟ�gG�ڕK�������K�j�(���P�0���Oe�}��D�����FR���� �`���5��j�ۭ��Q�5O;!Y����'�!)��m Qv�b�̋Do���ɀ��Tj���A��[�.�gԏ%R`	���sA��$���A��O�{ �=a�e�s��WLפ��3 F4���?�7|
��5 z�@' �������3�tQF�~��|N����oU�O�t��(�A �
6治�v�������TӜ��`�,b�FU���lk�z�G�vK������)����W�8Mrd���*�������:a�%������M�n4�N��X�/�����/`~��w�q�Ԑ���- �/uG��2�߯خ;�@��+k����)�m����0�r
������J�e*B|��|D�m����_eM	�P#���>�p��t��ay�����"헱{r_����?C�rV�b���'Zsv|v� ���t�6M���D����3b��>�/TZJk�H�����$]*����Ѭh>FY�N(w	$zGCm��m��Oj�(W�i�<c$*Ic{�(�c�mv�m�]���wWX��<�VQc �(S�V�T��W�n�YE�R��Y�%*�'���د�m����f�2�_�-�`���t���N~rܠ}T����*ASI�U�ǘ8��}+@˿�W6b�M*�"��Ih{B.���ڬDLI��4�86�T{�<W���>�iڕ�K�x� �d����Z�� ��l��XW�v&Z�N[�:M��&��}�L�_x�[_��z��Q�����u�Z���e��fWB�{�F\o!����]C�PJ��R������`������R��md���������[���~��f �٥z1z7E��E�k�]� ӥL�>�p��XŮ>ہc���@@fQg���1�u`�|k������6)"&؋:yOR��&�G4�Q�X�+��=�� �t��{�j8���,.O���Jy�I�-"%E�`�����OxߣCkXqE�<�띡���d+5�V�A�ں/?[�`o��Ϫ�}����/�R᬴��ԚՋa@���l]	,�_`��pS ;8��Ұ��?�Hc��խ���T%ȯ@
a����3:��T�f~!�SنA'�ɴ{k�3R��=��������(����Ƚj�䅵�!E4ܢ�?3k�;͟�rԟ�fF��.C�S6%�L�t33����-��/3,n�t\�[��o�|�MM����Fg���9�8����i�?a Rͩ��Xf^�J(���_�jYW p��@`��s��QTiLÖک����j�M^�;0�q8�7�[�G�(f�/��G1���A��C[��x����>��O)!8�!�cǿ/��.g�&KG�D�L-z%�N�l�����.f�,����0�﬘G�`(Q��
Ц�5�HD��F~�@F�E�Dl��5)�N��x��W1:�Y�_���e7������pO�W�BrW|##��>�3oT
K6:o��Dh45��ʀw����^-͌C�(�RB���\'P�<���9p#(�6udYg�c����@-�U�A6���������"6�b��'�<￼nZg�7�6i�SIvcc���� .tM2��1Z� �<�̽0.�4�۰��Zo�����zm-_ I'/>����xo�Z,Qvj�)���0No�8kI<���RVg�+a�1Uqz�ލ,���7�qz^�{�d��I,nM�fCr�1�KT�����r�|gu���C�~���y�F\�[�"H�����MJ���5�̯���ly��d���N��!Y�S��a�!�pEWJ���~���FȒv`�E-�Bb�凔?(����34K}��3ҨF�(�F���#�m=ri��g,z�c���KY?�YptXN��^��Wz�0��r�_	P�#=�3d���t�i�P��s:�	R���͸^	 ���T˧p(F�:���.h��Y+�|���
��� {lkmRp��U�T<���D�
�/�g��~�J�2�]��fo�#M5��%�z��VՆ� <��ʲ�k]�J�T�� �[�C_��!���~��y��c����r��{�����Tb��.]�m�$�f~1#��/O{A���0�
b�I`�:�n6��f��f�t}O#;i��gD�z�%�e�>q����z
3.�fs\�Ky�v�A=�C/�$�s�x�I�ɏA����\kNJ���W��UHWJm�CL��|08)g3~>-b~Rh� 0�eq4y4sGa�%��+���R�d�q��Dn6���F=��R��(g�wkf^?���Q��K�7��3	���cRK�.B��c���D�T�y48�3L��q��_V���[֣}%��y���IlΊ�nk��3�V=M=k��j{A�X�������;��9bn|���-���bmJ�r�8j�e��+ٍ��i���p�nֳ_��fwX�f�c;�:��زl<^ƺ����Zi��v��ѡ�)7h��F�!>,�r������&�d���ovϑ���(�,�"~Ma�u��+������߷��a�j\j��DHkfDr���<��y5q5{�\�� p�23љ\�v���y4�h�9j���޶9^�7P�ky4�ِP���	�͗�\~9��m�6�s�c�[@vn���I�p��H�������#��۵���0��f[N�?��6p�Xq��
@=�Ұ�x}��T��Kx�4�B5��Np�COo+��&ȟ�и���1���#��c�e��\(����v�e���HW�x���>Oc��[��b&1F�$ߜ����t1.����B��b�f����BqC&���(V#����d�aS�E�V��Ʊ�w����ү!ZD�x�"�)�F�O;W'/B�TT�at��rs�\7"�5t8�f(�����H<�_lĨc�' b���&pO���o̻M,�: ��Q�D��ݼ�#ˉ3����VS���&��LR�����s��=�.����Kk)�'��]�ᨉ��BaO2z`=�禆��5ԆwmWQ2�ߡw&�߇��|;"W}9a2t�
;`�2�^6W�T"��#������"rp|�
`H�P�в<n���l�K�@�ݹ���`hŊ���kL-�iVǠ��|oǰ�F,"ܸ��臷���l-�L���Xk����f�sL�3-{97��aT��_�,�+�q�ޥ��g㳍�F�fu��0[E��#
�x����yA�J��1�Rωَ���J�ѡkN|��+a���s(e������<�{�X�k�����]�es�M\�(�v��@�mHÏ!E��Jz�`
��*4�3�*�4L
�lB5���'�6�;2y�ゔE.�\�;IM&n߶"ѐ	 �Cjռ��)x���n�T�Op�_�B�	m���e�~�xUT��Ț���ި��Ҩ7��?(ڔ�i��9v������G���/T�޶6�*,LY��g��e@�+d��̎L��%��@�{}�#q�>5X�h��m5���2��Yi^ �MV#Tʬ��������D����� &��ls,��i�5����6o�u51+�J4�S8��#�G�UΈ1�mogG�E��(��YJ~{�҆+GO��oʸ�ЊmEAεQ���!�;
�<�IW�(�?ߕ/KC�X�V)�w	��0�oN]bX��6fd���qr^�]ԕ��y!f�f���R],�â�c�8�ƐJ��,���͘_�����&U�&}�"�*��H��2u[����h���y�Ҩ7����	-tj髦�R�ؤ"�I�av���(\!�7H�X
�~�������NAh�4��x���|6��dL=A�oJX����;5�i�v��Y�c���8|SZ�fm��w�_��!i�w�/\-��\v���h"
�~�������:|��o�w�O�M�{~��m]�{�<�N�O� �(��hX��v��3w��+�v\���y�nyLo�L]� ��Հ|I�Ϻ:I�?��3h���59�5�W=��\7��]O})s��.����4������t��.��
��DcF������T*�J��Ba�4eR�K���,.�ɕOs@$S�+j�
f���?nk�1�4�Ϙ^�t�A���c�C+>�S�Zc�v�2N���l"��Eď�>��`m��<�UMi1��G�r���[f�=	���c�$�G\���TX���h}H��j���R�|�r���5�㡱��J��` �1@�y��J$��
4��{)�Y��*�Ԝ0.�Ot��d����=�w37D4��}|��Z	;��#!�2�o͸��Il� �x�[#Ku�3�q��%S�� �KE(��^1>J;��\0�D�[�6D#����u{-|3fVx���99���w�*Ի�U���ʰn��w
R�{᜞P+���T�K��[|.��%���ϱk֐��?:�>����j���
���)u�F)e�#hJ~�Bqk�L��`>���_��_�Ѵ;s�����K0L�nE��raY��怠��@�a��vwIo0�Kl/�̃Ԧ.�-�i�U%�CL�wqF7@��Q
X�@;��A�\�\Z����ks�k��=����)X\�NT��} fJV��!	�Y�^%��*̗�J�-�&hAB�>ԥ�JW�ڀ�i����f��Nʕ���J8Р��a$��Nx{�x��Ԉl��?�^�ѮEjۜ�� ~�8�hǥ����,����-x��N�ѣdG������gߞ�_|���a~����&U���*����tl��x�J6�gh��+��N� 9>Cw%y�I���4��B0�YT�|y%la¾E��{�@.X�Ű�F�g]�g�:����ņM=�V�Ϩ�<iR��k��o��ϻdeWi�.��L���7��S����Y�;W��B�,��@NRp��ܝ�*���a�t/��,~���:%��_&��;Usu���FDP�x���ƪ%~C:0�j|�n+������u'.��r�^�a�U�&���im�nv�/�]T�U�{����׀�$�Gm(���� @�������
�^�`0�b�0s�m ��j��
s��-���?��8��������"=_
����,zG[�	^���Y�蠎���Mr�n�~��H�i����* ��uH&a�+�v5���.t�Y9,T����!��ݪ|�Vd869��5����2g�y�`7y�_ ��=<s!��SK�;<���Yj�e�Z���/ܕ,�����[��������[�vF�� opf��G��������Á7�K99q�8gP��}����Fɯ�<�/��7���/IȽ�<)N&�i
>)�*�#��� �����W�HLXgL���K���SNy�����)O�VǾ废Yo[��\av��$f���1>�ek"zIc�'qD'���]�a��2(�rk�>	��y��`��������Ԅlix�Mc��C���8�!lb"�Tsw���L�:q��Y�NԐ*�
sc8X]��O����^s#v.kp�<��Ϭ8#�n?'�[�SUd�+�����F8����.w
���w��I������!�%�O���'ʧ|7�%yY}o��>�$"ɩ�ru��������C�j���jg8�C���r����8��"�3n����VN���!2��Js%��%� ��-��nV��;9 �b��D}$3�8l�
�a���0ى��%����#yG�#_L!W���=t��	�f+X(H�)QA����DE�	q:��K�`�AZ��Zo�����{a.��m˥�ǧ_�楠�ú\Q����e��U�?��z{4(�$�l�,��y �qld��g����b��t�T����"%�2�O0%�<C��hi�����
9��#qK���C?I6��!Hӓ��)��=,G�f���O�K�N�	�dtH!�����b9��f�=s�>,-$�I)�s�c����өk��n�e�{�R��8��E��r�����g���:W璅��������)��s�v(|[*����|�Z%ξ�������wV**1.�"�w%��e���L���Ѣ  BalI�tW���3=Xq��J��(�4Q�V��G�[|T���w3�����<f�W�c}����^�Í��^�H(m':��H���ag��#Z�J��P�(�k�&*C`Ğ1��*��M�PH�[��Ȃ@\h��u��;O�	&��%�(�>ñ��pM�(B�bw���ľ� D=�H�
q�i��ZI0����,r��Bj�o
!h��p�$�aH�1���p##%�c3"l
^�d�I�D���?���+�&�^�/X?��%O蛝iOy�ol��l�4Y��ka�53�|��1@T�d�cm#K��J��\D$ u}�ʦ��ј�W _W�H���z�>��j1�k k�'w����R��Tl��F�k�%��������S���.Eű���@;w� ����[Yi^����\7,�Ѝ����&��O�jS��Ҋ���0��Jo����U����LĊ|6<:�* ��՗�����5ϕH�.R��k1�)��#5�����4�u2!��"�Xw�w�;�@��p�Ħ�\��R���5�p�B�˄<l�ҩ�f�u,.��x�C� �p�2A��l��J��۶,��g`�aғ<���R �J
{ Or/��C�O�@�7�j�Gl�O������L����~�`	}�{I�� ������I+=�)���k�K��l�BQ��<7 Z�@��],f���3e����RM��0�YS��n2��5����p�VF.�3B����a�u��Ve8!RC� uc,�f��]P��i���6�sJ�6���Z=�RM���ȀD<�F>�J���H�+��Q�s��ây�s1�%)�rafP��"꨾�u4=1}��c1`K�0��B©\���X�&���w���і\)b��5��:������8�p�0��u���@͜� B�{t,'�7ôw��*T/�#EK2�%��y�� ��%J���k��z���������/�zv�m�^r�afk�ڒ'r����aI���jE�Ε�j��j� 5 �5�	j
g�x˰܌�z_�����.?2_��Do=�^]����kA��i���l#�T���T@n�]��P���_�B�C�鶕7��
�.S��'I7��b'N�!ټK��R����,.�]z�z^%�>v�+���� rgWL��l=�M4�3��1�'��Mv#�z�_C�١�m�N�}�24Xﭏ��r���V�F���d�O�x�%��q�,%�jQ٠ؗU-H��V^�v�}~`�7�}�cV��M�aN�зA��qD�^2چ!�K#��F�E^��NmN}�U�U:t�	 �v�dww/��B_ㇿ�̵�����f
�I'O0h�m�x5h(tǥ��%�b�n%^ўH~!��N��[%�����*�*}��ͮ�D33<�K�_}�H-e��jetDq����My�D�ٛ�̚`~C��vgh�-+�1��j�f���Siӑ$*j4
V��b)kˏ��s��f}2\�gR ˹���G�b�Ws���"L�+�fg	��W�@1y�����]U�A�����hsڋ��{��C4*��얜�+�^ٽ�f;��_��M���%�WX��֎�uO��'�b�i?���7~3%6,_��s-?`^M�@̻�X�Na��~b&�
HJܝ�Aͯ��?�|��"z�
����x�����8�x U����X���~WX����@�^���=K.t���M���KlGK��C0	��r�¾zh���os�'���DT��F���D?�� @�8zw&͊�~�M�+wP�ĕ��pS�,���-pl�J�*�̵c�c�Y�$%l��bT	�8���kt�xړ%m\&p�M�o_��q� ��=Te� ���]H�#ʬ�YhX���h|�>�0��3%Cd�fJ����Ύ�D a�|�W��Vױ�g@�k�чi��k�p��ٓ$��M�C7����ML6;,%�(����a�5H>��������I� �	�"z��<0��E=� ��X �C!X-G�6��ܥV�3� ��i�K��y��/, K��וŊ��ØÔ~닶G\��hd�� m+k����-M���i�1� $^��wTP�iQ�g�ݒ�.s����v~�葔o�<������qʮ�t'��7�)L���4�%�FY)q�VĀ�I���bG�@�D����� G�6�������4ݟ�Rk��!Yg�+\	_�B��t��e�	Lv�V����4<�` �0��=�
����$E�I�q���\�����C$��r������h�Eև��5���Dn�>j�s1����4��_f�(V�]Q�)�dD�ݱs�C�Y��H`�#'�o�ij�N���B�	���K��U����1��rR,��� W����)�ʥ�M�W`m���A��Lஸ�2�gK��e�������հ*a�ϵ+"6��;\Oz�Ēvt�p�n���J����F�Y6X
�'{>���x~xZNV��B>[���WG�˾9��z�S`Y^FԮ���n�&ILh`�Ϗ��u�{��۹�����%���%g�V��-O>����~���G�^*[�[��M�K���#�4\�&�|<V��$�τ׊#j��w��C����+h����1�Z�}Q�
�G�Ke��,�9�9`��pX������*�VL�"�ł�8C�q6�����z�M �~$��	يܫ2�_���:�O�C0a�A̧�6�v�� ��x2�ùK_d�QB�B��z��"��v�:<f�F��,A��?�Η�㷣q��u�[�`$� M��,.��My.كz�`X���<�9E�Ǆ�.T_$�捣^7T�t�T&��C�/y���""f�D,���p���`�+0<�odH[+�\Ft.&=��!JP��>�13�
�V�r���������VMJ$�\��[��l(L��i?01hS�wZ47Q���4������P��W�w)�{KfXl)(r�y���r���$�-�09��u�:h ?���|���>$��S��!�YM����[�/�Z��ۚT��H<��n�Ɋ�*:���"��T��b��s�⺦%�N�Ρ�Dj�h!_���E\� �Y��=
�R�\ z�.c_�j;�������m�^10��<5�L�굤��9�հ|�CV�f+?.uNG�n�GB9���[�2�TmH��7���JVh��2�1h���'4�.\l�E�%c���ǫ��&�V��tt�Ǥ�
��9�}y���S̒�-},�Ce�^�*P���8Ǫ!ƹ��3o��:[�P��h�}���b��!���`.�%Vb)f��$�X����A��a�Y��펇�|&�-Jp�r=�H��I
O��7/�%�S{�#��i�>s��c��ҭ)1����K�m�I5�-��]�4x�ޑi��?��(��W>�_e��/�ܤ��-��hlf|�R�N��x�=���#�����G/B���ڨ�&:���m�����A���p�����]pr�j2��a�ĥ�L�D����Ǧˢt ς�9��sS�Df�	���� ��Z�$?�y�Fhl�oZ��A>"^#;����ޑ���[��c����0�֧���9�@^f�p)E�.��t��"#�:� BI:�;:�%\Wl�^�<ݘ�����6<�[�
,{�"(캦����l��q��܌qz����]�n>�?v�P63}�<���K���;(��餴0g��۶ß!^^�:+�]��4�BWqY{�'`f'�'���f�#�5	a��5��$�+Cf0�|4'.A.���_��ƅ�+�}ּh�c��������&/\W<֤�׻� %�/��{������^��|�m�|�EU�<V!�)�Ji�K����jeV)��������.#�:�b ��v^�P��b��M��Ĩ,�Ow�/��*��]4����A������Sᙈ�`��4m��{�7�J�k��V��Z�1��P���@�ZD2��O��;yN�gN@s��d��yV�#���_:Q�+�Ż�gPZ,]����GL�L�0R�^����bS:��nV�JwgB��j��^�q�`�p� ��@f���u?�q)Uafn���0��G��Dt���}�6�g��%��C�)f�����DЅ:ƨ���0QI+�G��
����%���aV�c�&:`*"`.�EU����f��_ɀ�r�t�6]#�gB���T�T��w�3?�4'F8�����㷐��e�X�o���n�����x�^����-`���tC�pw�GKMYN��9���k[l����y8�U��=~U.�:�V
5�~nj�E^Q��VSqJ�?��)���#������+��LZ&IN�("��	t��M�D�88�m��6�d(q������H�Oķ�5}x�r�E[�X#���['� ���|t�ERٍ��� ϼ[��/7��
ix���$��3p8�/��J���Z� ���d��l��7�7 �b�.q��jmT&#-�2��z����l[ة��,&Ū$*��A���4ܕ�ʹY#��^�P^^�#�[���hXr�F�^]��*+�S��4"��B�����r0g�7B�C��@��Q�~��׵gæȜ���|������H eCè�א+Pݞ�,�(l�e�]�b����M~��&��X�z�_��(C8`�䪣�	y�� �s[�k��nh���aW�l��o���(��/���㼮�aN���6������/�ʗS���{��/�I�r3�������6ja��
��g�&�ְ�z��G�����m��J�W����]��t��/��@�fW�b�/�N���������� w����XT�'��t�#u�KHt�����saɻ�妛� ��he��L6���A�!�Tч�i���fc-=��A�0.H~�4�o��M}�W���`Q�Ie ��%�49�rtaZ2F��0�)�P����2��C׏����������1��D�ђ��8��{�8^R�{�	���/�թ�e[���:k'�luV�D�'kV�c���[m��`�YZ�4%Y��	��#�R�+U`���|�S�Zu_+&��Ad\��{�A���}�Xj�l�V�#}��MC�<��������v��^��%���`�OL��^[�R����PJך��j�jg�_������?��\�C5[�m�:Q��q`~��O2:R.f����.�$���^���<�����cHr4d�]��܎춣�H���Ԍ���p	��	��a2���d�J̸ؾ��9B����	�)E�Ez� D��P[�L�l��=]�tX3��Nf0g�%��S�̇ ���7' �����T��7�.u�q|��Qi�e0qw<Z?���W��;�k�m]T�-F�����_�p)p����W���+dF.��;a��,�n�e�*1��y\{ѧ�\��[B���kb�dp�R^�-W�9>���h��pw��۔�S�aw���������PJ�&��/�����\�E6wвT}1Y
nt�e՟E.#�S���̡4̉�4*Cv���*�ŞL��˯�娆��z͈cy�ԁnA�NR�0>�%���r��kA���w���g	�+�P93Q�'��6_E����0G�(�}I��]�]pt��cx�����m&����]hwt�OA�6�� �f"��!��w����ofc��r����q�Ζ��R�C[>��;W2�����C�+�A��h��߶����r7���GyN�)o�N�6�"�D!��\� �H���k�լ\���eD|��S�!:�oI�O�4@�!M!x粿���KJ??�F�U��~])D���A�}��!�Q���V�~��7�>�`�N�|g��#{~�- �̽xC?㊤|��{�M��g���<��p��� z�nw�GT:ļ�!�mp#�yN	5�YDa܇(,��"߀�6x�3��И��)�FSo���\���v%1�QL�͒��������o���4�3+�=�����r����5"�i�IWS����Lׂ2G���S�����x��LTp��yOç���G�|���]�	��1'\sZp?#p"qŠS<�^1��d����wy]k��ひJ�d5�'N�'nT�^ZG�xdp)�|���P\�y�����ފ�q�O0u(Ȇ/1�Na�}��!�'V��A7@��$��At�6r�U%���/}��r������`���" ~�c��b�2d�%GP;�r��`C�_3���pU��/enu��R��q�u�=��ʓ�-�1��O�Kfs�Rd��Q,*�$�,�@ָ�R]a���\�ބݥ P�0"��;�N��#��á5\>t+nP���܄�9�R
-����/���A,��Vi�q���>B/3�����#x��$'P�ճd��z�Db����I��#{��x=N�
�&c�[�����I\�d����^Ӧ`~Ӄ���U��,=;�sv�F�Rg��G����j	�� -O.8Nc�y�������Q��'o�`�UT����ؓ�8	N��^֍���d��{[�"��Gsn�=ŧ��w2�.�Zr�k�@���'h�E���'\�&�$��la`Y!��#�{I�U��x�iS\��
%,�Kn]�Yj�a%eo����=p��Ҵ}.Wd�C��~�^(�@���=j��f�[{�]�W/ւx��~�ы�Z��'A�=�{�)s�����u&i��K�|8�~ڋ�O�nPt$! �^�E������Q7ҷb�� ���FBZ5�n��Y,\�'�x� g-�E�Y�v��^��T��YX�x2<�-���Z���Vk�𚫴��l�Vk�Y}O~v���-v-N�$U*��o�RBz�aO�O ��C�昆ː�~�B�Ph}S[��d@��AW��g	�wj�����uXXoE���D�4���0}���Z
��xDH;�v�Q��0S���M3�°��}x�m~��A��8�`q��.�6�	=�'�O���@X1��F����N^�����y֞��N�t0���b�ܟ���xhեm�}>��P��5�r�`�لؓ�e�#�z��g2�z��&��Q�j�c�2�:��D�G�	�#֭���N���8ލ���G`���������E����7��b�w)g55w��_�����Y6$�V�8���X��L�@�&��f�J��׽�M�o߹��4�w���1��˧F�4�n�B��Gm�������J��5�W�ANbW��T�u��F�����3J�2�6\�����t��nU%?��A�Etsb�޴�2m�vh�|�/KN�Q�2%\��zju!�<��B������f��~ƫ��E"l�[�+l�(,���0�`���t�@�c�<
��A�Y��B}7*�_4-���d��i��-|��\}��@��@��+�[0�,W�����5h���r�Nƽ������<��tN�L��J°��;<�����!"�6h�b)ؠ�.{C|�(�$Qѻe/��^�,���(_s�B�RW�[�h���!�k����V"�`�F]ћ�e:������ݧS�M|9N'���X�|[;z�G}ֳ���R-���=�'��'�w\�]N�Dċ��"$*�#���3��P����uA�����E^RDkR&�ݼ9�KK_��[��i��2�]�"k�|��m���c�{w���,9 �Ӑ�25�!��݌��ȣ6 	� \C[��6�tk.�~�t��fE��M�f�D#'�B#�emԣ���MSH�&��2�A�z�j��|����A����|3�����3���jY��H���ąN��n�+"m��9�9˃eW�KR�$K�1$Z���j�;~bdۢ��W�\"`8�P��ۆ�������� ���H5��R��G�Q3ټj���8rQ�p"0@q?Kc\U�h��Le�!f9�#�0R��ף�W�f�Y�H+Z;SO��cͪ�`.N����sgG���鏟t�" =��{���F�Sʯ�i����+]k@ǵ���G*�@�p�⋕l�pSl��_MQ�u�z:791��5km��u_��4��jH�\����%;E�+�%'I�ls9�<>�M�h�b�(�x�x����NB�i5d�ig5��х��%ľ�̍���aJ"�3�{@÷X��ի��v:dd�d'�ڹ���c�ʚ��4J_�F�L���!���m�WԹNiLxe,l���(pyA� }�@�m��i��jC�X��8¼������gՑ����^��?�h:x�n�kd�f �?D?�����DM��+Ɍ\. ��%޷Q8݁��ՙ��HD���4����aTg���k#��瘸C��E�9aA���Tq\=�[�`c��8lWr_b��@��b-����oƅ�d�H�t����}��)ڱ��U�e��@S?��V��[*Z�x��52��jl���`d!68-�dm׆�ђ�m�4Y�K<\\�Z#�읁%x�G%��tKX�.n��Q�C�O~o%/W�v�,����d��X/����w�~0޼M��l׺�!&l���Y���Kbã�)���L�n��_�Z� .�!�U�1�7x��Yy��J;�m��Z���Ҡ:z:[��b�j���~j�<v�0�����^q]�`�߼l(��A�N���c�����~�MY��Q�M4�$ȟ&%��Tp*K�^�_U|��W��;M��̃#Ì�%�l�En��;Y��J�⡹u�qMo���REA1ăl�
@�Ge�dWd<k_c	��n����u��
���>�lz��"%�4n�Kb1	.c�Z)������[��y-�?�¦s	��������Sś�tjc��(�܀���6��i���g��.$z�F�)�ydI��<��9Ƶ�L�X<a} P6�M55ƺ���a�E&�g��륮U�gxD�MӴ�ZE�ۊ
vޢ�x�_h���R�	�+�����9~���T �}I��.�jv��p���:<�^M�&q���[ދ��>4��']T���)���M{6�k��xI��ubC+�Ա�!U���&�w��]�-`V�
Y(y�&"ZB��}A��2ٮ���!H]�P!<�������"��\�q��[���|\�.x&��$���=_f[��	�	b����<��[��..��=G�ޣ�s�F��� c"��s��g�١#%�t݈NۄS.�p�%.�q ͷ2}�^<fj-�u��33��i���*j��^�����3Fo��cl�����AP���x�S��;Z��j�^�I���]��s��^#�
	$W�fu<�aռlu�ꡞ����ze�����T7�/V"�~l�+a�.�`sOQ�%����_1��4�[aG-*d]��Ȟ������Q�ƨ�f�z�DX�=2� Nm	D�n&퐸@Y�Bu	M��a�ұ�Cҥޅ��mn{X�Iv)) �B-��*��y4�M� ��F��.)Aa�D;T8V���2�jN� #rFo���XRk�'�
�d"!S�pI ���`�$~L��|p8�aUL���02�C�|���r�hp<}��c���mf�6/�&e�i����=w9Ĵݺ8B-�T,��ִ�ڰ�V��b��h��0d��5%�	71Dn��$,/�y3r��(���Y����m'd�N	u�F��V$@�VY�Y�3�_Z���mZ��<j.�^Gq�k�jz�#�c���ԵĎ������� �l�g�G����8���TB��Ҍ�9Ǝh�.:����0f�#6�fp�hyĴ���v�it�O�c8J��?ЮS�'L�W�w�?gA����Ơq�3ݿ�q���G�>Ie��u�ҕ�2��D69�8Tk���zVz�8v�u�jG���� ���Bx^�X����"QXH��v�T����<�jŴl�j�K��I�ג��!Թ_YW_��,�-�1��4������B��&#���4�0��j.6���"�x*��	/k��X�""�w/�5%��?{5WPn��ޑ]Xl��|mG%���?Ż�Ws��:��"��$�_r���<�*e]���ʥtD�Z�*Z�ʦ��O�1���Y5pa���M���`���=[���T�����Zt���Yo�=���r�����U��-�E�&��HF�y��F��^��>X�h���x�9G>�
,ޢ��(�a���w~��Dd�s��^ĝY�P�?k%qV���{󑍗�]�,����j�]��1u)i'I��I��.�O<8`JD��!�Շ��dq���8F���݉T4"a���}��Kbk�sHpPFа�ɮ��ŉF)Ķ�=V\��kB5�c+|���mf�6LzV�E��Qcҷ���n-M����Dug�b�MYz7ss�/*3�mLz�xS����B^߹�R:��Xi�a��F��ܗ1�p����:G'����R~Ҷ�6�<e�x4Kp�y�HL?D�tқ���?�V����+-ԝY�s�����	���=���1p$�o� >|~U$�G����Ux���R۾�
Ha~H���+K3ȕ�����B���ǉ�8G��}��;9���A��m��"�FӐ����ha��y��^(�i�[qQ3iu�b�}��0�lߌ��
�g�����X5�+e=����ּj
z@��3�u-`](�[�����,k�����o��Z^��q1���\�H�8�5i�m�pk�v��g��916��7gȋ����f���rxv1vb|��{"�[�baV00�35��C`.ԣ2g���GK7�Т%�5����H��մy����~����V������U��n�h�F����oK�q�U|p*��  �捽j�4!��,�X�t1Awsa�5
ޫv�,�Z���K{{_H'��6IN��d�`s�&FQ_���J���"�df&�A�0��yK��k(o��|h��m<xBr: }L�OT�a��J@_���)��w .��2�g�(�%�����[�9S�nR-eV�_���:L�\+��}�LE��4�1}C%��$�Œ�{����E-s��@���}�ƵI�����G�����B�g:���!�
�dG�a����SW�o��p�]5b�k�|�j��:�4�ݥ�y;�I|��1�n�j{͡%"r�=��>U�n}=�������8�nO9脮%�
�	�����n�[E�c͋�=�Ä@�[aC�/��G{m���s�DD]i*����>`�����.�9ɀ���̵��3����� ]#MmX ��s�pU���+�N�i�Y���dT�ó�8wYH/�`�/
H�;{m)s�Tf�yW���*��$��4�杍��	g7Y�<O[��=vL���9�B������*R�E �f	��<&\����I��5�K9�M��A9k�av�=�N�َ$S<��/���q��J�my�pGB��Ϧ�>R��K�O�F�#ebP��<��@2H>)�a�!	U�#q;/#mZ�X$Yd>n���%���6lɐspH�T�W��{��9�����H�"�h/(Fn����NֽS��p�=X�,t��>����k���N�eqxI��"�����w�M�"�̯|MW�-��Qx�����=��U��ï�0ցQ��}�d��r���p�����Xf��Yd��1���v�T�lV4mƘ�D��{�K$�]��BD��`Mʢ�r��W`<���Ĳ�x_�f�:ڜ��1)ݶ�u�{Q�羽����|�zZ���b8���1���Z�X?[4_�o���xG�Tr@E��c'��j��]��V��Y��ӭ<zY��RƄ�o�q��3n�z�%���t�fS`����`k3o'��0NS�SV��u�L��	���"�A0H����!�P�/��Id�\����t#�ؖȃ�q�G"���ĝ�A�LB�:���]�!�˅�����B<t�!�/�>�{�3 '���v�r;��A�,��b��N��E��T�;�[1��A^�ȸ�����đa���^�K�
ɴ��_F!
!De�� �m./4���-��ok���vF��F�>UșD]�H�α���������?�v���A��3�?�E��,M�f�Z�=���'3�N*"p&ZD�nE��"�� ���r"���l>���������c�E��}ׁ�c		P����!]P����y�3W�|{.A:�QPz�)[/�����bGc����zAG
<�>mq�YaA��u�N�.Ib�4N�+22���OkY�k.˷�=4�.��?��9�5�v;���dϘBv]��Y�A$�P��������)%
�FQlD��_ *�-#�9�[��I04��d�&�Bo�\��=��T���w�Z�b��~T�B�����?���mu�	f����i:��zZ4���J��y�r��L�Fڝ������HK [����:��A��uQ��^��K�7��h�(l�4���CeD��"�-���ʮ�}İ�~6Z���e5h��;B���|��b��Tz�?H�c7	�>o�К7�6�?f	H��x��b��n���,S/��a�����5�����'���BO[Κso�;v>' a�&<<Or��;2;O kNޜw�# �V��#kH�Iu�}Js# B��0��͎���U�9E$L���b{/�<��/qJ��q�٤J��Ĵ�x���q1F@�,/�����b���q���w��L�D?ZmB5+�@�N��R�՟�To��L���^"��,�BC�����>�R�=-��a�&�6>�}3��mޡD+x�TK��b���%K��@�/l��F�J�f�M��{��h��C![���)?��#��9�/`0�H㐽�M'��ĉ����;�pP6�O��O��O=;���ޒ��+���D�I���N(]��Y�����H6q0�g>(��Ձ�q��<?��>[y��ŵ
Υ�		U��C}������F̖puwO��Jb=�%�?�K����I��ܴ1q�6Ґ�L��<�Gز�� f,B�1� ��s+Z����8�f�_B>	�I*��{��*�}�Y�DQC�y��a�ɦ�_hy���7��l�^��6c[e�V�C��2c�w���Ez��K	�)��=D����YL?Hq��)�!�k��L6;}P*[�'R�Q�'�9��Xp`������P��u,��۵���[�ܩq�<��ߊÔ�X���qj�qHv���b`mPϨsM�d�?�d�p���V�?�%}�~Y!xա�w;�����������������%B���L�E�rț�cQ��V��h"�A�8:ksb떰��Wߢ_�s���o�K��؅��8Q���K�O�=@�g���Q��q����,�k���Ĵ&��Zg�j���&��-RgH<��_[��l��� ���A
��%b��MW��RQٹ1kN��0�c��.��v��e��*90(�҄"��?Z��.��O�g�<�|=�v�pYC�0z�Ƹ�֋p�?r�P�_gy���Vw��?=�R��� ڙ��n�Ft�XE7q��O��_>���A�d�#p��/\�Nt�?������6��E����X<O�O_�M��	�	A��b�(��z���M0޿�y�D����Ԭ�U�1�H*׬E���g�w���u�ɘ����z
s���9R��,����3H�t@����\7�f�o Sn�2|v)=���N�HB"Z�? �g"&h�WkH��rn��{l�`�ʖj�zos�.�<���e�O����e�bG�S��)|}z�0P��7�u�yi+�_:�"b��^A��T���[�Z�c��`��T�2�� 8皽X���F�`�ۉu��-��
��`X� ��	z�T�.4|0�}�a��<h/';|��7H��K�p��	�N����9u�Mc�@��aG��Z��6���'�&��d�f����*�T�_�Ч,����� t�F�
���:�"�7D��5h1^��hk�� � ��f�i��$�m���!�fm�`�ct��.Ǚ��-8Lǅ�	�ֽ]Y�O7��_j")VIE��e<�]��=�f���,�ي*��?�X}�Z���m��� a�1&��`����
6�1V	���e�KH�5* mM#XWq����.��x���VY�5���2�>M6�=HSO��>�6o0�t:��5+������m�8h�Q��E�@�]�cKOk/�u�V�s��7��N���l��T�I��/�aVd�B�u=��G�v0�9��L�4��V��"������2��9���pB�����;�* ��*��?���Ƒ�e�K�G~=��1�.Aݷ��0ӕ��֮�b�[�হ��:�<�P��ǿY둌���-E䝤��ލ��(g>-?����j�3�ʡ���T-ћ�8�|�4r��5�[um�.�`�}�8�5ܶ�@a�?��|�D�6�O2@w����MΫ�D�%cZ^� ��� j�:kq��>�2XZ� �Z����1�22�+HL5ח��P����Ӈ	6��m���Xd���uo�)��rX2��T��g��� �-x\x���V�B��AW�F�5n���zUч ���$-_qBl�q=�3ERotXu<�c\_��H4'��P�2ͮV��
,	014�ͩ�S�]�����
�a��	�ȁ��l���i>'�D����Z��n��a�އ��,k�3>�yȳ���9�®C�n�{��wc����������^��<��@�������3+��8��� (@�DL�k)�~�N���I�,&$����9���i�-��m�&�.,�	w�ȁ잴���WP�T]�ũM�R[�Ph�W���0zu��R�OWY��3Hx�ne����|�hC�Y��H�k��D��>ks��e�^�d��E&ޯ[���X��!�_�5t踦���3��8��@݅�u�)Ւ�d������"7J���6i�z�F�#��=ǯo�;nڰB�RZo��͇�Ӥ��z�ˠeb��GM�����j����/��(�l�_z��=�|F\L94C8Z�O��l�ȁ8w�wq���T�Y�F��e�����L�hn�2Y���wU�ݸ<!:�� h�;��^�j��� )��&��Z���V�:#W�ʜ��E���W��|�X���g���8�A��]",+l$�|����^bb�S[�Gz������ސ3W���I�yOɮ\`v�b>�V�ňF0{����>�0�!�:{�!l"G��"n�S��⋌�<#/W�p{�Q�\���l�4�����k/[�O��:S�	�=^�@�����SOεSVӕh�sT�M��<�G�vST;ڴޏJ%5�tC��nΦ��0�vx��A�Ȕ�N%M�7&�����QWl�sg�<�s��\ZL8�'kqHO��5������6��C �j$:�K��;Fy73�b�~�$Y4_�� ����|#����*����}:,%�b��,ʻW��̛��{��|�q�+�Q�OA�!�:Q�-���	LV�@B�&^>Pg`�	"�K��J]'[<RκI����o�ak<���3rߤœ�RQ�Ʋ��]�9�������Q�<�����N[�)�[�u��y��i�U,r�p�@m��7b!u���شZ<_vE!�(��ʩT�f�cZE�0`9�a�#"�@����_3��Z*Ɉ��ԮD�jDK@��6A�)y�+�\>y��m��Ћ&��+���2�"�@+M��5����/ψ�g/yax��$*M�Y �`�5�Z�Z�:�.`	z�'H�o�Bh�����g�OK��Z���#��x(s�<Rg��{��p�����x��
���H[�8��Uӂ��Wnu�u�9C�BR���a?���<I�S\z?��^�W3C2���������ޅW���F^�W���5?��`KkW�ޅm�έ-;Sz�t���-c�~�g��g>���|(��#5�.D�ɒ����a�����y���������&�-M��� ��c���Ry3 ��,��@46����0D������,�u������B � SoC�����I�C�ۑ$o%=�m�W-��q�7j�*��&p��]�ץo�sτ���YvB�:�:�f�����#k�P1��f�Z�V!�����e]TȀhm�2ɧ���U}Q�ăY�Dt���^ӰG�^y�ΖY���#�A�z�D�����u��K1(?6�����A;􅧼[Y��sڹ�dR�A�Jd3A9/�w0$d�h���9���c����f@?���tq8�z��Pd�#]�����������R<n�îc�9�3~7]���ȷ�<���4U�t:FN�ސs6�c	��}���p�c��vvǎ'���eȋgB��=(�rO-��$�\I�Gx�a@�E���:��L�zT!�����V���yר���Px�_�$��k�Cd��GO����^�\���t蟉�U���[q_9�}��ߍ��t��FC��3�H��[X-���`��zz�T{:����0�mE9�2��K��3���S"�>SM®V�hlŃb!��?o���7����
�A
*cq����X��g��dg�dn��^Z���.�q@�F[����n�1q�������nUeh	 �Xo@a�������������|���T�� �/�'.L��[���_2[�MK�����i���W����pE��Z��a����>I���Ti�m1a�Ԙ�I}Z�)��������n�ڤ�� �ۨ{�RU(��յ������:6��q٦��H����wd��S�p��^��VO ��P�m�</*�luH���`xZL��S�sf�"��f�}�m�2�_���N �С�G��ӟw��gXʃ:@s>��1���?xԫ�*j����z>��ϒg�Ӕ�pG���iBy�ʩ�]2_�n1e�t���<��gOn��c��=ר>�L�P��9F"�]srMc�e�c�Pp����NQD�"����I|@�F����X���7�8e���7k�3�vA�?����9U�����Ke8%��:�b]&4���<v�2:��h��F�K�e���!7�7�T�L�98&��(�-B[�1&ӨiWM���,�)G�i��R��y�B=�4ъY���m$DX8��I�&�Ł�S�A%��%.�.]�S����_����'ZdL�?0��;j����;��U9I�����a���I!�ܓawך��]Tde�����&��\�dc�d* a&�P�,�U�-f�DS�� W�g����уw�Ba�L��J%	�gR_���R���ݦK���}
7�
P�kg�v���03�2x��\�J��f�f�.V�)o�����|���>����'�_̇Z�FWCux�ƺ���3�]����`
&�����7B@���-4�Hӻ�a�C롇��Hij�KF����W?��0��Y�%-���)_ <��3��]��� h�
�Cc|J^Pq���Ht�ɨ�2*}�,g�i.�=]u�_y��gdr�c�v�	�.F�xT`{T.-��Dq烪���V��f���2ݑ�<�ta;��T����;X�Zr��f""�{�9�~/�h�B�`3j��l�%C{�qN�I Z0���I��
G�`-�_&��*ED����KS�?�rrѓ����'�Ȧ�
I8��i�t�b��c�V	��ꘫ����8�K�a�eM�Q7n�ȓ�Dt���s��'��׻,�^A��&���w� �� %T<^�Һ�����Ps�q��j�?���*
ٗ.ach�qC[�L+W�@i����Պ�d��z$?T�5�5 ��V۸�>����E�mO�!S{��c?"sf0F���WzH�(��!��d*iҰ.�R�����]G�S>wH�`<�}`��Y<-
|�eWq�R^c��}4a�����\)o���>��_��C��z�"/��T�����ɦ�7E�~�>����I�qf9h��(��SS֗�}RL�J�턵
/�����'�l%��2��z^�P��ot�Ef�N7 &�}чY���	�k榻
�grz����u�~�I�����pT�E�]���J��[3>��?捧�Ҧ���������g��{()�	���a�KH����."t)d���pE���1��:�D��+��EH4��� m���x�YI�Y˻��x'�8,�o8��:�N�rG@#�i���O%ʄ{琽�H�qo�翚tA%ќ}�>�X�B߷���8:���)��7
�)����jX�ɣ��~u�ѳ ��,�;�@VV����Xf`(��ZjV#S�9A��e	Ѕt@N�,jS�^�Ո�,-����;��2��:6��(e������C05:�����o��Z�5eW��T~L�u?��ɞ��~@6�Ut��^4 �m�������]'�h�A�	5�� �e����e���$Z1w5��SA�j�:0/�w-��!f	��9��l�ۉ� 
��/�8�1�B*n_t�S�]�g�U�����%�ΤK>{8��կ�R�35��=#��>�ښUo(K����u�w�A�Wuh;?� �H�����~$Qn	��%���Ҿ7�3�{�q�wv1�%��sJ��Hz����!�*Gzo�����Q�FĬ���K�A`���l�8��TPg�v]�������/��2]���߉�8��'3�>SՈ�P$�O��k�H���ÇM�f�/b[Bg$^r��x.%��HgFڂ3m!��׎�O�X���b���4�zJ�7X��$�r���.�9�{����vy�̗ ϻ
p
Ld/q���*�M����	�A,c�J�fͮd��h����sw�|[&�0�<�	k��(�#"��Ԟ5y|�d� ��	ΘDjSe�2W���KOE5�����Leg0yH@��L;��e����]�������T��=k�j�̗%���7����<`ܢ{�O���.sJݹ6���_;��82K�ť/}�ȯ��i����~lD��\�p�YC�`�fgT�`��a�ۓ��3�9����5�`Hb���{Gf{q�_j=���˳'T��`��dZ��qY���-n[.ka�3�u���A]�="�{�˲qv�ZyU��^���R� ���D
9n����7��:إB�9����G?-�/aÝB�L��JJ۟&������ڹR�??;e4���pPs���?����Ԋɤ��*��/�h�����ヵ�0��u���o:�qk�&��}[օ� #sB�FJ�(Nf���"S��<�� ֧��3~ҏ��o�niU���OE�6򏕟������ǰ�!� <vc�iY���)�;94�we����٦zR�?9�@��i.�`/w�%p�sV]{�1���կX���u�/�vh��-��\���N�b<7&�� a����z̫�I�h��FX�w�1��]"�4W�凍+�^�6�E��]�A">̼����R�G��~^m����}�]��_d8�����Q1ܻ�c��Ը���$'ה����)pd1��	A�О��BR�Q������lm��Q�F�ֿ�,+����pGf{��lƇ/���$�|Ӷ,{����D���UX�&A�0���k�[0�	��Q6�7|[Dɞ�@Ș9w�i�T3�,�?��ݛ�P��81�~Ε�f��FK�ݽu�=�����x嶿o ���-��t���7�͐o�%L8HӸ��] #��lGFC"�?+��)7ɖ{깼�P�|M㉝�z@~�K߁�L����7u^Я��)u97�h+��'ܥ>�Pn���"�.��*'^I�8Ү�0A�Z�0��W�˥Ԙ2�
��t�H�Q����u��3��h�l�8�g�E�`�Vի�L`�ai���#�F)?��~�ܸH��gu�h���S�)9�R��<h��C4��,�O��5����ᪿ"H�6�ֹ���r`�{_t8���{�<��d����[������ʒV�ՒO��U��c�Z��m�q�3U�Ӛ�(�#;�1K��Nl@���
ϋ�ʔ�(��O7���f0�RI���ջH{0��ۘQ��3���E�/������	�E"�a�K-dd)gr��s�RpqV����P7�Ȣ��j�W�c�([>wL��셸u��&6�c2�\?��S	}�C�a'�Zh����WJe�����W��&>�K�� &U$�'���ٹT��	ܱ���Tt;J"ԏ��+{���V�uT�>�rz�Iwœ3yC7�O4d*\�OTm��S4��f����A[+~Q
$q(h�xJ-��G���K.;t߄��	}$'���*h)������&w�)�����,��|~�ew�C��d܉�r2�k�cnmP�����x��y���#a?�쐢����=7lh%]G���ڕ�*u'�x�U6H�*������"�J`�b4j.s��wE%[��&����pgv�w���b��{KG0yד��R�Q�愱OZ�kW�B��يa�/��^]���k�LnY([�TG8/VDh�E(>:����DU`Xl������ �����/�l�U��Pm�A�^��g��m�1)�,g��Q׌��yn��g:E�#cW������g͉Q�(+���&g�ZB��W���g������|��k����O5�-�@�/�-�A҇(���xb��qb�ѝ��3QH��=��(@��&�J�+��S��?���~�i=�pL��R���G��r�ouo�(6�d�u3uyt2{_��E��n�?�a����C���/��nL��fz�l�I
�.�^=��RU���Z����b��H.�I3��(a���Ҵ�fhJ�4 �ZF���t/\ 5h�0�_�NZ����shW�Vs��փk��qk*jΑ�`>����щ�߀.��z�E?+5�}�������;���q�&�I�+\��R{�H�=wV� t�*��{H]�Z_���Іx3~�s'�3���}��/fr��B��t���t֒�P?�ho���\,�2���M�2x�="BU�gT��+4��֦`�3OF$AX+� ��$��2���y�o�gb�]Hi�'{��B;�j�F�����u�	x��L�m�D�(q�v�.����D�C��j�1z��Z8@QpU]2� .��=ac+$��Q6����GN�f{K�	�	��`u@�h(Qt���-j*߈p��$13D��eQA�4t3�^XCin��'���(r��}�?�c�Lx�h�Ѽ�@���nly("��M���;���$�T��#��]��~b�ɦ�!x����kb�v��Q�������W�57f��="����砆������I;�T�7m�E�܀>�ͽ8���x����j������q♄�����^�'��k�����ob�}�ܵl�bP\���&�z���E=�w�ם(�J�B�}�зp�����Cl�5��
j�ڣ�z�Ҍ7�s����2��U%�^z��/��A�%G+�C���\�sk���+tAp\�ڮ�	�Sa�OA,#5���*,$b����ZA�3�+(�����b���"A�ԡ%��r��S5 �4�0q�g]�"_	*Uqs?�Ke��V��7]�R)�#p|�,6�H�rRt�萋�cy�b֞ �#���`�Eh�|���h] ���l]	Z��|���p�,���Fļ�P�ڮ���3 �!����Rf�x+H%�X\/�a峅���t=>ߖ7p]�� �Н�M���#y5���� �A ���=��Y�oе�^q,�C���m#ĭ�J�j"v��7iq)��0/F&W���n�uI
�V0�S����_Y��	`�q�v�1�I{���W[����~˶:§�tK ��ì�}!r'�fn&��b����9{���[1���U:��T���_��Z7]����"������;�_������� _YJ�/f��*��<;!����=��F\&����إb-�-Nw�ӊ���S]Ҍ�i� ��M��*P�.u&Y�����ܒ�v}���,9��&t|�]�F�fŴ�{JGje$������;���'-�(�t遳.-��d�Eס���~5
T�:OO��!���v]����((���K�vj�My�x	$
�a���Q{#������-v���Z�'��3�>IOߘ<��Pԙw�OM��Y���"����F�i�ˬ}���p6��؃�%�#.��$�w|c��6�VM6��~
�!«h�S�����:�������J��^᮸��k�N��*�\�Y�
F�M�����a�� ��$�{)�]/Dw� �O͕OS;����Y��Z1��欗���45�F�Y�=��o�]VKZ`W�B��&] j���;�֎�03�/������F�%�	�1�I���6�9�XqN��ǳ1������
D�B�E��HPB�9��P���:��R�"��0W/
��w�Ǳ�-M��ఊ|���S�7�����U�Ci˷�Q�/��4�����]Y�^�\Ѽu�qxr�4�f�:L,+�&�ּ�!8Lb6�>`��_�tUD�;J|�LV�j�H!��`2�d��yC^�0\��-�NGJF<��<'jC�n`�V����E+��2ekZ��!�tB���ul"~_g}X�m�:���(�T��!�h��������h�� n^2�,��ߏ/�/�ɮT���~��Z����]��3
���qA�*�k�֑0h�fV-o6��DP����M���Y�s�JcSx�^���������	 i4�4|B̛X�;M�B���cv�;W�����P�q_�]So��6��Z�
�Ż7�\�&.7�8`8:Q��],�T����?�N^�w%���$���-7ц�	�n��V ��r8X������Ҫ��e���	����NЙ��i�u]dJ�'%�X2!��*Ъ ���i�ͤ*����~i����%{����ƺ^��q�C,ӘFS>T�Θ֥"���^��K����">�e�q�h�'��P�D��^]8���o:����/�n��=aΪ�=�=�f�zC����Z���HqF�]�b����TQ���iAR�=(H�l��	��ò|�1�ݡ��3Ȅt�N˵��2��LN���7b�ņ{��[��sz��x�)�AP�K܂�Ɍ:D2gY��ħKT
����e�AMF[��-��@��@K��4V�o��7]-n^+@:H?)}�a��~�+�%z�:��5��%�X����{Xn6ɷl'C�Ĩ��p+D�R+�8̧� $͍�M1�PyŶb
Ш�id�|CX��G	z��i;�'�{cHi����G'`�<'�P��m�$��=T�S�1��v2���
�����!�( > BYC1�X&ɔ��C�

)�%��H(H�lnN\ތ�$�&(Cc0\`<��������W��12`�s��=Ho��Z�ދ�� ��6���D��Đ�w�Md�Wd��z���� �M:~u�3S���ATJ7u��of�y�41�8�F�sM&�K��WNB�{<Tg[�F���Y�#iw�`'|ص�>�Y\ɾ� ��s�~v�d��kib���:|K��OYg�ސ�U���S������0��-+�T"��j�g�E�z�<�v�� C�א��A7� �B�ń�5�>�i��S�!o�E�2!�PE7�φ��s���/��U��D��g[{d7�	%u��6A�
�jL�Р{	b�J�n�S̺S����m�����Ē��!���PL�*XW�n;nq�M���~1{M}$��chi��)���%^-�#M�Fܧ�ÇBuRA>u�I�N�F%E7�'P��ƩkB�]���l�C
���6)��rTTL��_TR��yd�D��bGC{}���u��<�P�8D���!9��x���-U�Kؠ��]_]� ?�)c&��_3�N��4�S��	��*�wydϡ�ye�ӿ~[�Մ����bʎl��k{��{Z��|���(wd����ݣ��Ak�;�
3y�K����< vم��!Ɇ�
���~���]r�K,$OWjc����7q��7���2�o�K��̸C�6@�8�4��#�#/�&��s /xd�Ŧ$��&&����YC�]IS63k�O��p�`@�H�(�J���de�SK�+�z%�x�hܳL~yl�Ay�P��`B܃p��긯���ɰ�m%��cQ�G����HH�aJog��?�w�D}�0G�\ɽ<e��k��I#�*Vf�D���4P�)w	/����{��4��]Z����i؁�><G�����M�Jo�`�CuY�\���ҝ�������B���A� ��LRKd"�fY�FQoW��|1.��&K̏����D�*���2���t������toם�	Gm�)Z��Q���!
d.Ѵ+X(�U
��e��'�hd�E�Zޱ7�����`�^�I7ː&�ο(EI�2�_�`aR��e-�.]����4�[��KU����˞�.��4�q1�|����B'�k՗{Q�*����ƞ���H�~6��P����,�@�v��a�[P�6�4c�p����c	��өi#x�!���d*;z�զ��<Іv�5-~�bv�K4�|��M���)n���o��ߗ�k�ۄu������-0�\�h	�'T*a�#qgU���w���bCJl�I�0�'Bj���f����sqܰu���(t��V �U�[���¤���Q�a�9`z��u)��:�N.� ��v�QV���Y��.����-��Ck�)�]�*D���(���ws=�b2�{��#��b^��E,h����Ar@��
�ݑ/�@."�t{٥��p/����Qvi���8�
	������� ���C��
�Z/`('�J�d�CQ������}����1�2��q>O�b�r���#��Qkmf5�b��O����ޕqfC����Ӗ�(O���+��ւ�������I�Q�O�4��kΉ�QƐ��$�I��L^�ɂ�4}���͆e�)Y���ccS����W��*�RW`��Ȳ�_٥~����"��a!%V�/�������(ܿC�a�^�<��]�+�j���S���B���%��ׁԕ�z����u��u�yL-�9'�٢�i�Do�{�.����~֖������D���dU�-L���y9�k:I0h���y����*犘ںY��C��d�
y�T4�<�i�������R�H{g!�a~
j^d-�m��eYo����EN��Go"�5�NF�lp�AJ�d���v�ൂ�����ȍ�	���&��&��)�c���e�� �š�c���ڼ�[��w���B"Dq�0˜���T�A�����TE{i\{2^�4X�+���7܋f#�k�3F��N�����>V��E��hG�Bdm��X*(I��*t�߃xx�E�.=ˢ}��V�4hc9�/���s�����-b���/�����b�cŜ/�2����96A�h?��#��d%l���H߄J'ѣ�{�������
 $g�W���o��xk�ޝ���,���i.il�,������mk��fB�
���`�!A\��'���x�l��I?���f�� \n�'�@���8�wlI��*XՋ�^���\T�୦��F V�j���m,o͛t%��HH<��.�{�l���2�(�J�8<��9~��EWC�#ܔ���(J�4�>����In���
�gg��g��x$�������̨�D��EsK�gk���;�"���`��P^�����+����<����a_�daU��4L�F��hy����%M0 �:��ν4�o���b<7��xk�kXh����F�R�i�N*H�vID)w�4�xУ��L�r��f����_�WQ����P����)$D��X܇q�xL�x��԰�}ܦdb��h����7e���.[j�|X.��iDVW�'W���G1����%O���J(���ҋ벑�?ꖻ���C�Hn�V���=g���K����T4ֽ�p �N�Hp���kinX�޾ղ�I�ˡEo?GkQ��R��W�!��� O�A���vB�U�@X�v��s�$rD6/��bn��G��<�p�qX�'	��Vlx�ꕆ� m�ۺ\Ȥ1�~0[{�Ѷ�O�:�p�c_�����7H��L-P�e	�z!�r�����M����	w��[���j�5ȘO�?ŏ�v�/��ɦ�ߜ�ؾp�|pz}��4���kN����!��@	����yR�,�����g���
��BK2�zu��X*W;����Q���F���ꇙ&,�j���J3F�{��������z��+d��"ɛc�C!��)��BՔp9�0虵�u5�@b����So�;�E�&]�;��s�����VcH*Aӭ��*o��6�����7��N<R^e����l��=�F1@c�ۯ���xagW������y�'Pk� ����d���U�m�2�M��M�^���
#���?���G%�l�G���tf8����V��+�P'�x,�<�8�e�M&��;A�U��z�Ie�	�2�2��7Q��hT6?��?��WE��1[8|�z[���Ƨ�5�}(ª2�XVo���3C��f���U�b��8��L���8+k��:s�Nt�H�Ь�)�%3֤�S�.@sh۲BJkE��>�5$� �����$�M��B��߱S0Xu�I� H��w���H�r�V�D8wP��
uǖM��\E���v�^���-���[�\S�G���=���qy��V�Ȟ�;)`o\��N@�������QmՂ.���a�������o�o�w����COTp]�ð��i4awq	y+�(G���qIR2�4��P"��t^R�<B�cc��aԣe0�+��e�6\�����oH⶟�Q��'��rb��;��7z��t�0k~���H�i�?s]*�l�)Fq�o�§�Se��_�Ol�ൂ'w�$���G��@$N��;<[\d���j�U�e�Gb�`�S=?�[~����i���֞�?-�eGI���Y�I�ߌ�_n?q�9�6��!��،��(�S��~,&�nLoQ�\�Vi�dG�\���'�I�	NC=��)������z�p�M8�u�oz$�~5���qpT�Y7�$�{@��T���u�)���/��(�u�Dey��&�	�O0�K�lo��1��$����߽����������Ix�m�,y���=A��Y���*Ŋk��q���#Z�� �^�e6;��%�*��0{�0�*��!r@s��S�$:���O�@'����7M;�w����~��wG�����-���ԗ������R�������3��;�¦����)���z1F����3�q�3�J(���8;����2~� �r9|�'���8�F�j�y��d��]&6T�6!�P�W��C�c�G���_ܥ�g�]�_��E�Q�f�YW��Ǖl�mVMW���=���--�ғ��Zf[2��:&�[t�M9�8Z�HC�S7?��*2>�gG~�R�_�>f9�4�D��y�lU]jN�:2Nzz���Ċ�{
M��<�=��8�W�$�xl�1W�d1c����zy��Ρ���Hı��m�t!?�� �!��f�P���R�����d}�M|.�E����ZRX��;{�6��~sȜ!{��@� �����-����Շ}�w�&l�����k��dJ�`b"֣�#���!��Y��'ƪiX���({�h9|K�(���T)�4��_�͋�~+������Q��T&i�ro?0�~=�П9�:�nU	qAt���T�I���ζ����ƾ��#���,>א�n@�
��$�"6CbJ����\�E}l�.�1��,�Y�M�В��%RƲ��b{ά�h�����n��R"nd�!0�����G`(U�O��q-�8@�^l���L�z�e;@pΜwV,�-��p�Q�	�vK|$��
"gҠgm�w
���x.G�ؒ�Y#�#�����k�����p$�Ep��n��_�s	Ʌ��lTʧo�kgGW�@��w��5������jl��h7wD���%��9��,������󿆻��wH��BK��dN?Z���J�%�9#?���g߭�9n�HX�>?wKw�+?
����4l���vO�@��4S���FI�tYG
`����26��ӵn�l�s�L�d�#b|����j�.�Z�& �|=;��/�,w��qx�:3����g�<����tT��٨ػ�a�9"\ ��EX��^Uao$>���N�\.̖א��.����3��˙���p~WM�����>�ȏ�n$�ҝzv�<��ܟI9ɧ�*� �b5$x�%�����;$�b�D���:�c5�:��4�c�`��޽ڽ��T�SMz��D�+o��04Q��ZJ�����S����|_@�p�jr�z�+<N8���-�iVme��FP�ˇ����VD'n�q:C�1(������7�Qu�����I�̇�:)M��k5L�n��e+���}�o~Ϟ(o�L���8��L �L֕d���ׅ�����<��+,[��;��Mp9̒^��f�q�Rf�s�')qٯ��y�X?4�S�+?,R+Wt�s�����d��s�y�V���N� ��F)�>��3�J��+���>��(��}\�q�I	w�?�C8ҫJ���
^�v�k�M�n�F߭g�uZ$o��md�f���1�Ɏ�ԣ�&��Nl�
e��V(�������*<-�~O����bE4�ѠB�~d�g���Sn�%`�-~G��4���r���/�.l��}Yb�3x�♨!��5���Y��a�^��ؒt��ϴ2J|ߕ6���D/pP?��b���-L�B�R��r1ؗ�[����O�n��\f��]���'�� i�CV`?�N�X��
��>w�Us��U�}�n��-���	�� 1�A�Q8�z9	(�cj�{�x×ql!1��L5st2`�fl-f4�l�����;�e�DQe���νjLّ�i�b�e���|�a�z΋�-�R��BV������Е�"ʎv�H�+&q�6_���F�!�Z
+4f>�6	�!q�ˑ,q�`����������Rζ���ܓ#]v����m���#aJ��¦*�,��^�|C��n��P��g�8����0L�	,(,�j���:%���w�l���@)�0��3��/���p]�h���D���u
4uK7�Q�qL�M���[úa����v�⨭�zI�{��+V|�C3��������ʭ,�W�8 %k�W+#f��)�l��N>з������b���z���?�@G�������\h4~�H�Ay�{N��Cӎo�S�����u�Ε(:�3�僈��2�[eL�]�b{ �}�t���W7(IkEU�Rt���I�8�wf�4�g#tEK�<m* ;=t��*�^���=��k�C�jމ�RjNgs(�My��xRu:�r��} �ǒ��9�2�5���{?l��4�լ�g�DQ���I��@;Y�n�	��H�1�������-�|p���1�N��}��y��lx5��������{mvb���-(����X��ߙmk&�ܔ��76�ɷW�CX�Zc�J��� R���+o�$�G?V��&<� ��434h�F!��;��V���+-WF�U
�E�>e/�,��<��k�W��E�w�$��F
�P����ߒ��k,B�����Ӕ9Ni@X�0��L`�>�[�K��F/<v�mSr�k�����t7���{X�g>#��r襖/⊯07��t�!9ʊ(�^
)y&�-���%������\b��M<�H�� �h��}�h0.>K`��_��	�}f��nW�r��yFF���S��*��W��Lb^�q�H�H=�U�8~v����9�U�YG,:c�t��0�g���P���	�z�?���	��2�
�O����bл�K9'�t�Jv�E�u�y�$�����%�w{��|g+��� �i=*&m����#S[�()�/U�@�B�Y��
$2�S�`=Q"!)�� ȍ/o~��5�2��Ʀ���R��shl��r-)����K�h���m@�A ��+-4�U�uin#NR!g������̉�U�֓�#���_��h���û�C�'�`	��L���Ni_���O�p;�iط�[��\�|i򰍉���rC0/wtğjg�;Q��D,������as��Ɖ�ɉh,��q�rP��0�:�Ύ������2����g��x�DJf$;7���-�
��q�V�WC�ǵ)N	��̪�R��Z|��p���gX@on�s	��懾���v����uT�-fqP�B�I�G��1(�¨��қ�ɔ�f,�_p�Q-�;Qƫ/�>����/Z�wK������s�>IL�ȂT3�/����9 ��˷���|� �>��(KmJ�� ��̟��n�h��0j�:��$�#a�n
"�H�KpT����0s��/�5X�Ke��V�WUtԬ�]���`�㱫7>�-���Oz��G�������0Y�;�.�������>>r���O�Vt�j�cAb�>��Jao����X5�U�v���2dD�QKb�hZ'V]5G�����B�n}J��V-��aj��v���p���@�?(H���p��"2ߴ��p#U,y�� �C�$�c�o#p��g��b�cQER�Z+�_���1@5��m�����U��w���oUF���jF�@Z�n*��NV��ײ�{�/��(),�U=�J�����ޞ0�t��o��aR:؞h(h��yx�#eg���47(V�93i��OD�� �_HN��BCD�ep���τ&��&�EZ���hC/�A�U�H�NL��̝�N�INS��h�cY]�)�&,��N�Yi=@o��ɔL��|=8�킲o{�����\!ۥ�X�m�pb���E�G)�#{ڦ'�� �!�;�1����*�a�YD��$+��YdƁj�/8��:�S�@.B��A�JG&�s��)RHQ��#$��Hy��t�|{�Ρ�qʔ�� "S�\)����&�H�D�仢��{��ߨ��a=�*����<�XN+���t�D�W��5�ՎJ �c�5
��D���pM�2r�k���б�Ht$���<��!���*��5&1ACaR����>C՝T8��h�����\]:�OK��2���/vP�4���܍��i%�b���g����*���R��܃n��}��`^[�R
��R�?�G?n��p�S��L��W���hR�� ���S���oxL�DfR��=��׈K���T8$fʠ�g91pG��͏mm� ��R "��N�k��,v�@S,�=B���������?��8ό��>�(z+Ovk�2Q^���Q-��j`�T}yo�I�ӟf)��B��x!���![<|�؈Z���jcϖ�A���+"��
ɞ�
�V��W��E���-�Jh�Ϲ�s�@��ǿ�kq��M6�Dw���O(�Vj+�]��y7+&Z�=�Tv��p�s����0x"�ͣe_�J�0'j-����Y���h�3S1���#�{\YEU�Hp�qc�x�[57�϶�]ٕ�p�6a1S&���{?/��R�ً���2�H�m��*��)�Hͨ����
�k�וG��b^���"�q���gi;xw�v[��)Ǔp[[\茳�|�,g,��P�j���Uҟ�V�.�~��>9�Ws�zA,��CS� (A��� �/|\�dM�`w{N�Gv�W�p���k)��ҟ���H�s��7$̌SN��*�c�~�+��ԁ0�a����	9�#��hc�p�w��� B�ң��J?�=8�~���v�2���i֚#��%�L���N!J{�B3R�Ȏ�����D�^~�&L���v�[8�Q&:r(Я�'o<#�̕g�OQ��k��nI��m{I6�DF�:MR���������z�����+�!(ީ��ܡ��@���S�Jf�H�Cu:�Z�owx�#�{<,L�E�"�|�Z�V�}�Ǹww�{-���
p��j�H+�]���N�TS�f���W2XR��Йc����uwe�Í���k�tFDT):�Ϭ�Ƴt��1����΍e�L��Y��.詗3CR���n�7dS~ �:������Ѿg�X.\�4��RV2�ZqtI�N��Ȟq���>[�c�l���I�3F��+�ᩍ$p-:"��Nuk���W�]��>8���b;m�޷���c_�UiF�ǐ"���6oXA�|���17@�qM��Лӱ�R��J$E������&�qbW��� "�{\�(4MNp�8�6|��^R�
����g�)���@�x���q�� �������Ϯ��)A���7x���}��u�b�������z3̱,��� �Pci6��沖VP��Qu���[��0iNB��T�(��T��������{:C��{Yd;�;;)����%Ҏ�?��`4n��m�S07����N_��;�%�p׳|du�V���;=6뻰I&n�q(!���n�%���R�����vR&�{�fi<���-~�!�Nj}dX��|=��c�V���L�H|f�w�z��T��mމS�����&�j��T���b|�̖l������]�.�d����rHP "/{�6��_��GN[K�gL�m������O;��]�߉p�R��fi�@E�1�,��K���Z��&Kl��%�ৣ�C���S%�9 ���`�4a���M��^U�>��n��S�*�c�hc���1N|X�-�t7�І��	�)��T���b R�Ü��o�[���,�!Ђrm�SO���0O_?�P|U�����{>�W�:�Q�:��T����	���i<�-�({��p6Fq��E��, p:W�r����Z|Z�xL�+M�yV������c�&�aŸ�)?	C0��Q$���.忪;��8�P,��l�G���ٷ=CB]:S�>���tew�(��!�e�^r���dtCU��]�Uj�2y��MM��dǃ�����L��S�Q���f�� ���f�'r�����［��~��~��I�p,	�i���TN���[�%ً��L�*��`:Ǫ��W�lV�����֝�����R|�I+F�
��^��A�����PNy���7[�]&}b}n3ذB]�-�P��qm����-J����U-���� Qc�?�������4��#@F����qh��|���K}��{�4�T�&&E�F���j)M�[�s�/���x,�`6x�e�yo��`)V]P*����1s����N��\&�X�@a���F��鈐�Oo�{�FU�+��9Ǳn����HH4f�0�@W�DU�)���t���](E��[<����[< .�~�l���tX�QgҔ��r}B��}d�W�����VlrV���H d�9�eN�~3��9�x�/�e��OC�ܘ&�{�k��H]H~q=~DJ�M�P"P��۩$�,�IB���\xȫ�E�VC�����@H5�q{�H����[���.�EEkM�2m�_���61�J{���Z=��UW�]��Adע���]$�w�a���x����xoEUQ��N ��ruquڍw瘰�U��8w�>����J�zm��6�����0?�>�VK��^m2�z*bc����,J�C���Z��𶬱�ϛr�#ξ����Ԓ�@���`B�e��P0Ld�%P$�I-�{zC��k�Ҡ�՝�R�\�6�8[�
� M��\�xp����S���,[J�Wy��lG�`Z�JGį��c�LoC�.~N��|�X���|��?�C�uM��(���uWż�&��~�ಮf����BqS�Ғ{�� ����a0�B�6w|��o��H{��P�!b��N�=��I�}���q�:�b�6(���?ϩK��3����.�%Q����_��5\<����aJ��}�r�N�s=���Z�}�S9�V&܆���C��ꛮ*�n1l�u�j"(J�15=�z�KS���WeAi	N���r���:���4V���e.F��w���|��iY�&}�������b�.���^�i�X� Ɠ��)��^C{��9i�ל��HZl�H�TS��1��>��V����p}^��'njۨON��+�h�Ar����>m{t��^yp�N�	`�qE�f�m��>���u��XT͂�%,3���>>�I![܁ߥZ+��}r`�pt������"6��X" �^b�e̸������z+�XBc%٥"~�����޺9�PV}a��<��&������R9��������],��1Β�1�pf��%̎ p�}� �%��0��0���s�Βpj�����4���D�Kl���/U��%��ui��Ga�;n�c�l�:���x�Nrf���~.��c�5l�Q%+�_L� ��.1[3hH`��QP,7b�Y�r��u���e�DS��������i��8�D\���f�')��vf���ҋ�Zj0�
S~�C�ps��u��*���5k?�vFR{/+�Z����U��L�?�����;���	ZA?�U�L��ѝA��,��85��^=&4���uBw�!�71�L��r�f�n��B�}��8��='O}�5gGd^-�7��[׬8�3�^V~��d���;�J�b8C��?�>��p�ȓrY��a��G�/���oy�t�3�O�Tf�1��GA�'��O0��7��>*)�2��<�"�2`=�O�_�l��Y���c�m�)�+x3,��F��X���GՄ=l�$������x/|���q����c�t6�/6>��fP@�6�f�!�v��$�#�1��+qK�m�����y%���A�t�CАVu w�� *��A"Қ���.= g���d����4y���_[|��U�-�ꯋ��@�{� �p�K���f��7����i/Es+"�-SN`de[;#1B�f=���^����=�9cأ��[��i�;�����[}��,�
�W��5)��*''�s8�<M`iU`�*n��@�6,�-�
������z½K����r�$NpKph�gz���H�N�ėsǙ�i��͘��P�Y�;� �Sua�r��v�7`�QB(�5X��fm�J_L%�]���\�݀�t�+/ǁ5�� �Z�Ё\F7�B�+�G�鷇I!S+����cA�����c3�@��E���`udT88�X�����_M���[AQJ��՚�0'Ƚw��-pg�����h��v��5tO̳�\�<.�K��-�Gر$.
'��}~��3��+A�$��Ҳs���Ql���۪�4�u�LҺU�����i����c)��)�ة�l8w~�3m����Lş_Wn��橵%����t���~"]�y��KG���s���x��f|�����ڻ�c�bZ��-���&�n��N�m�k)ʅ[���Y}��I:dU��ܮ!�M��J3߹ֲv�N9��P�MN�8ޖ�;洛zf�st)��gN��w�%���;�G�䴈�C����@��BE�`�"QP�'a��Qh#N�N�Z�c�	��3/Zm*��6��,�Y�
������*�E^��s��6�Z4��k$�ȭ����)��I͙�K�Os�A*�1*�.[�8`/+�0����1ٝ�wj6��8R�ǅ�p�wy��TSk��Wľ1��ޅur��(��ѥ�;���"�y�9	���5��q�~�f"��A����+^���O�zE��	��c���:�S�P�����Ҏ0h�F��J����~.fK&��+e=���/#i}�ǒ�'�6x=ڱf�'E��̥�.144*�,#���?� J_M�4��DV��Џ��g�LQ�D{
l^`@煆��&�s�
�b���O�W�:�"h�熈c��LH���7�ޑ@���Ž5��N\�
��u#�Sq�4Gʛ���}E7�W�P�`e��6��lP��x��x'K��;���ZRT��%�^�y��a�O�p@\����Τh���a���Յ`��?���L��i�:lD�[A�ʄ������&��U���[�6 xDIbM*����oJ��x_����k�^[u�@�_��q�hh�CV�����6���J��5�&W��V�
�e�5ڋ�"��5]�c�
@�W��J��L2zS,�K{�&K{�A�ȋ	1�	״e�)����!�&T��[��
)�����ٰ��L؝���M�툩T�>%��I�|�F��Yd`��TV+ʅ\�Ȋʢ�G9i%��-���??B~{�fQ�<�h�6���,~�!�%@=r�F�0f�U�]��K2�]�W���iK����X�#Ri(��.���L�>�^��������e���>ښ�\�z�+=�$�l"K���2�#��D�%���!)Q�A��9��|L��
�y�ai���f�E��Ϻ�SF8�aC���7�z�a���������r��,�%����[lYL�����_����v�~"iX��"dצ�d��s��;eK���2�.���n0$��IҾX�z��瓬N����8/7p�ω�R2�:xĮEt+���:��_�.T]\1��E�z�t����A	�4l�DȠx�p�/6���Q&c��:��a�	�]~��x�|���L�L�H६C�D�d	r��К%U�M�X�(❁5+�nh�#��b`�(T+��-�C�&Hs�';8ݾks�1l4�x��D�h��ʂ,�[��� 6]�.T�^�U��w\*�\�.in�����vtf�EC�U��o~��m�X��@�'�yY�S4���y��፲P�����V���b���'��rD��}����6�=�n�9҆�*�����o�!9\n3oUT��a@�iKJ���@�y��X$1#�%�@���B�Y"R�R���b��y9���΍�E�X'�9�CJ٤�I���|3�9�!�l�?)bo�������9���`� {A*�Y�u�>7.����C�*�WF�y �t���E�Mu�0��{I��h���Xrv� �F-��a��l7-�$���(}����?_N�/�*y_r��y�b��Mis�Ի\���o�!�?F��W�7�H�#��|~������=�/��6��(?{�[��8K�\U��m&Pv�ްQ��`�|z,�0��lj�m8���������<E��	t�Ж��|Dȏ~�c���V�t�w[`���1fG��'���S%<5-j�܋��J.�L�!NsJ1��� �� ~��H�OWP���m��L�����4JK�ԛ3Q�턲�`�X����(T�B�y���(��}j��r�d's�B�v�Q�����~�������nP�bgy���l�3aO�fQ�$}�j)*B���, +�E����E��Z�r��+��H䓤zk�{�ײ��3�f	�Y~�!�$|���!k���}�5�s��|��˂a'Ss��-��-bb�ή����n
�L��i���˲�;"��ΨE?�ɯ9йK�i�'�'��{ZA"Khϗ�4T���;uMv���6;��o�=t�
� U;/��g)$K�Tk+/�f�n�H�����axqWc�z��,����ң�ǯHIJʱ)�;�b�Z��r�(Ո��d/sU��|���{�_#���c~Z?-���^^�K)Ԃ�6-�[�6��|k}	�S�
�'�������W�X��i.�_�����(qd�^I�g�B!��-�d���$����G҃At6
o)�u�_����vy೨�n=3�I~��I��>ص9�����Ы;��xN�b1ϰ���ϥ���d9�{2~wׯ���LkM��U~��"�m	��9����Ӧ� F.@�c���Q���u���ey�J�����fRH_�ɯ�a��}"��$��t�x�}�ZN��u�c7۽h5�Y@�K���iQ%�^$����c�BZ5�N��OG�䔐�|�`c��"� GyZX�=��=�a.0[�
[:d�|�]$���h!�/@{�/Z�Ѳvl7�}���!�lT܎�Ch�g%��B��٨�`.X;v�v�)G뤩����Z��r"�ҥԗ�܆?'��G����nq<2�v/\$�&Wom��Yv���:��ጚ��g���
/{>81� �|,�,�@��ā�h�ō�����UU0�]x6ř�dV��D�[�I���0M��6�E��)T+Ȩ&�G�V\Jo%�V@���l�g�G���m�(����+D��Q�ѿ0�9����	1��KpK\�1G�!�Y!֊������Q]PC�&Ϫ�v#�ڲ�iU#�點��#t�3jWR�9��/Op���bX�Pwm��i�~�@`�2�#\a��-.���xA���� a�j|<��B�`B�)��Q�;��ly�XgF�%`�j�6�,aR�}�j�cM0�rJaA
Nc�&_��S����Fz��:��!B����N�����w�g���	�w0���\h�7�$��v{�a�f�=	���ak��.{�
wߵ�xf�'d�x�Ƣ@F%iU�p�X�RHl�\.=��@�l�%���u�gro,3��"�ԟ}��n%���>�</M�%��go��&�x$o���]�~T�#�`_�Z31��� �㶨������f-���HNe��ƘǐE?1t�����e���Z�����k0�W�sSi���D�Z^�P��htT�8}R�kD�8�ߒq=Q@yI��A�������o�.�"�b�)G^~�0�#�2)�}��1 ��D"	���E�֑YD�9K#1�T�&e��JO��An����J2�2N]ؼ�}�k~���I���g�<89�T	�:`�~^�HX�h{y��۸�d}{���*�cH��\��4e�
�o8�S!x�y�?e]���o�xc{ߐ�@	�"��Π��쭄���Dp��tb8�$)M����Ѽn���z,�
I�!5`ƥ�T����X{�a&!˓�7,��:�-��������°��,�,pn@G`_��z��o�&gbKT..=����������lst&�М�"����WW
�@��������"����J��� K��8m��_�Z՝�!%r�/Պ�x3� ~�oADh���l�!$D�ڥJO�w��GY\d��]�r�ir_U�5�x��9&�}��$?�m�9r����տ�����I�{��]�w��L��)Z_���X�i@�G1/f����n.	9@���FܺE�ݬr���n��l�`ͮ8*U��qP�e�W5!��k�m�e�ǔ߭�!R\��%�jr���⣺��M����\��^f�0P)9���-Ԙ�T��>��-��ne��gU;d4nzԂ�����/���o�W0u��H�/J�p�O�߄#�d�y���u}
$':�1c%q�� W6���+���g!��9��V!�T�Z���yf���^����k���" ֪3�F_$o9���#^������1����^8�����G�)��v��_ǟ�k><�J���mg%��n޽yf�#�z@[2>x
&D��#!Ɛ"���|�A�Q$fꪶV9թ�X�)�W=Vf{�T6��&�9���L�	l���g�:���e�b�0Ժ��%M�r��d�3r���II�����S��w(]o�~��h�@nTl��]<� �z2�2��,i>��(|ʔ��ﵢ����.�n1myn_$*�څ)2yJ#����Xz����B�+�(M��<p++�16`��GꇍJ˲����n��\�.���~�z�4/��U�n"�����ֈ�������ݠ�yg�D�X]� ��:ĆБ���~�70e~ؔ>#��}?xH���$�hs�d:q 4�a��x�,���3��i׾
�'M������m�u��܉��3�0yI$��·���k��h+0��
v���;��?��V�K9��y��S�������|��4s�lҝ	{�X1в7� � Q�aF��DMO�E��C~�ɤ�*��k�NE�Px�34/Є~�L�[t���ބwT��W[w�m����m�)���h�o�E�%�><-��N�����ȶ4g������B;�	&�x�p����]?Օ�F�"��?C5��/[���:����@�:��b��M�NȷFA��Z�.� 	��rUh˵DZ����Ԯ�-��M"������-}�ǩ�����Q�,�<f�����d�H��_�@όZ���tk˱f:s�Pݢ�;�7�3�)e��^��>��l��z6M�ш�n��u~�Z��3�|us`���C~��}��5�b�������g�Ike�*��}B���C���B� 	�(�l�^���Ԅ�B>��)�H/�Ƚ��Ԑ�/�:V}�ZýU
�U	�~g+g�F-��_���l$�N.{:ߠb���Si穥܆ҡ�O��C��<��X���k�|��ܝ}��ɵ�T�$뻆W� �I��<B0WK�?r_z�PI�wX����u�h�G������m��B80��޵�i��xM-�M��C����]�;Ϡ�&m �N�+��}C�z��i,Ղ~�U=����um�� x� ��ĞL�;�
"<�G3q��>�>9b����B���Q50�l����Xf�I�8����#�]Cr�!-D� W��n���+�.��f3{��i��=�V�,�l��`Z�V�.y��X�>�4�+H���ݝ����?H�A@f��6朷n���jD�P�t,`�m�6gHI��O�q��MR�X��<��F�&(P���V�]�թɉB��� :p{맒O_�D�m,Qt}�S��'����J�4�j�5�t{����q�ˣv��4�0*	���<rILd�D><��\���gz�QȗqmTT�g"�$�p�#Ճ;Q��k5)�R�d���<��o�ϗ�d�9���Mh�Ln��#�q$fcZѕ�MV���VeM����x�I����R����Y���'�h�ꥀ��F����?��ʟ��&��$�v?�TDϽ5��*�u�N��[*�~bں�g�!/֒-�B���@G�T(�L4�,�n�4�����/1��|�f�����z�2[GI冈���	`&������������K��ly�6�ȣrF�¡�ѽq�8Mp[ ��&�M�� �&i0������|�c���E�ի��}a��"eh�`I��:�[}��1�Y��|/���k]�X�r15��p�n3�]m?������B@X�����e+�����⤖��0�X���.^]����C}�=^�}E����~��@�9�;v�j{����������gF���;:��/=��v0U�Ow��t-y�T��]�#%��YT�ӗ�����j$�X.g"�����*�9�/�J
IC�R�2[*;�^y�"��Z}>1�7]��xF��"a�܇���K~��;(�A� 0�=�wG< d��W�%*+���f_�_�G�����1sv�;�����h�C���x�_���_=�f9�M�l�Ea3"�hEGfa���.`�"_��gt)j��C�6�G��d<:�x�m� W�N��w�v���6���m�e���u�ّ0Fdz�h�P�x�_m� ֱ�'��"ow�X�)�M���<�|̀�st����xO?"R���_��C|��A��$�I�$}���;�Sꗐ�ԡ�� 	�m^��/�˛"����glg��z�.}$3�ش��p6O�R�H�y��X*�T��0��I��!N���u��S�%��ꪗ�� �m���]����2vDP5���<,pZ{0��/�� �O�Ǡ�o=��D��|fja���]۬ڗ����yv�D��U�k6?�Z�֙W+K��}��C��-,@YT���DJ���JV�0���k�r�2Z�WhfC�\=��ڷ0&���(FSt��DWI��uN8�r�tШL�G�y�;���j~F� G�Ӵ�o�
�t�������p3�����Dj��)�]�-}�#l~q�=�� !�~7�a;Ѭ���LX��Q�<��_ƴ��
�6��;�<\�a�
^��g,�~�a�-�-��*2i"�K�)p430c1}-$ܹs!�0���rt�~��YLD���q�БM�Sӯ}�I��{� NJ{t�<D��%������H9kuO"wW�aq�j��5[�V�"��*g)����E�ْd{ink�rm�~�9I-$�X�"qф%�CsI8I{i������R(@�Q�f��{IwN�?�����M��ke�����!d%�A�Ի�	�S_��)�U�O�6���|<���z/0�����z���P��-�?�B�|��d����2V�L!�lI��" ���g�3�������^>�#�BF�<@���D�$ED�}�?�d�Rsn�6b�VXR�R�#yRw�ƕPˬԼ���P�2��ɋ�2k�ҩy��D;4^<�Cc�X�5��[A�r�bS��|�!�c�V7��$�r�8��2{���G��X&��*��=���-!w�*�O?5x\qn_l��y���Plu{3��nq��^����P������V�,In]#�m��L���7K��{��D��gIG�v�z���F�J�M������Ttu�k�!��"���1x�ק/��Oũ�E�T3.����^��_��_�o��w>�U ���6�(~� \~[U��h���e�h����E��cFE�i�w��G(�y�3��_���`���˱�¾!�]7~OA��Z�;������U���*d�1_�-ͻF4����nd�nUtœ�ϩ��W��-�/�`-y K}�k�����9��ǿ�	����� �8�O��j<�^7�#[�#�]�GX�KXj�+iOk��7+SV�<H:O�CH��PTqs�@A�dCn���<*���w�ѸUА!T��I�q�WX����i����)�΋o���=D���q���|?�>�v�0���\qi�!�ʼkyUo?��)*^��xj
�qџ��`����E��=9��l��9<)�Ӵ7QP����ɑ�����jDi;�-v7�B=�6��Rg���\r���@J�4��k�b�nض�,�H�ɠ�3���as��?B���2Rk,��1X�!�u��/�R2W�)�hc�R]��4��U/J�u㍧l�ǐ;��c|	�p�k���Eb�;��/����A� @!bf���;|'S� �,�lu4����Nd�E
�7��E:6�Y�V�aF�a
rvC�~�v�ӛ��+Kf2#S��fXx���EYG���e��^�uR%Q���q����Y~:Ϙ.mR�7t��_�.��ř��:���-5��hl#a��a ��h�/C��Ln�����-�NΡԺ��� ǔh���_¿<��[�S-�mP�ɔ$���}(�x�R1�X���QB�M5��f/�e���E�:��"��'#�\YC�9�77t�)��7ws_�>#��^?Z<�Ĭ>b`$`McK8��Q��<n�.�O������z�?��l�1EO�P��,ؽ�ϖ�.�z�[ �ޯ*�9�"8��t|��p7�w3,\���s�y�?P|�'��\bPr�K�x�n�i�b��p�%\�:��(���JfZ�|�J�W�t���'i��	��R6ٌ��?>����g~�˪�h��SF�	U�6�T�k��Qt�k�W8�7$��2�h�%&]��Y�'$WvA��y������K�懲M�]ب���T�V���,���1��`�
w�Q�*y���(��-B�y�P�}�07b_I��=��V!���9%x�A���l^f�M�g�f6Tm�Rݦ���j���r��u�0��sZ�'�KQt�	e6*����,�n��	��������2!r2�1N19P�guZC;��;H��ዑ�cd#�B��kd��U�;���G�� ����_��ꍇ�{��U� ן�/��oC�������L�p�����e�G�?�.O7�������!e�1���Qc�V�/�P�!(ܠ�< ۦE�3��x[����ߒ�K����!���#��c��)�(I�]�y��ј_���Q�3g��Un}c	:B��i	��⾰F6�n�^V�9G��|��]�q8�f䧦�&hЁ�U�?� w�!÷�E�N��:�}l��{x�9tU�5��MLL=7R���Y������+�oy�� � �o���>�;+"��LgO?䜱��q2{�P����sWfh��(3J�L���X�y!���QZs(�Q��]E����S�i���V��բ!^F��_:��]�V�V#Xԙ�<��ɮx� ����D����离B2�=�F��!��M��)M��Rɰ�=y�������A|&^�
Z��w���|�&�<P�cW�Y~+��:o�dL��`�)��|Yl~��>Sp��qX����5��uDf	�15P�y�s���m}a��(�l}*��桾�:����$GN{�W��hK/�ށ�P�kp������B��v����,�B�X~�E u����������~���i���'2!&p%B���{x� ��b�n͢Q�����V���~���`3%a����H�X��K���.!�VG��a-�j�A?Ă�����F!�ʂ��1[� ��h�ݒ������Ǩ9=�jSۙ�|iT��h$�^-�:��� HS�:�6TR�$H��7f�#��vp�& E'��<�|xgnK�{/�9���*�j�NA�f������4���a�!ze���J��gEW��Z�v�-Ti��������B���&$��"rC�a�0㓡���e��@>V�|�AFH���oԀ������W�������$e>��I��\�qtAL�_2�S]E 
P����Z�Ƌ�ð�Iin-*Z�GE3����F��er�!\����J_�%	o�4i����Q����	A�gW���g�-�Q I��V�U�Թ��Y�;��v����u斬,���Qt,�(Eѥع�\lv��]|�$"4��^�1B���X8>zBĭM?�U��J��W�\��N5�6|�����ٔ����.@�D-�`���'�uL�p�/U7*$ٓ6'U˜�}�}֔i���ŤUa/�x��&q����OK�2�N9���A#fpy�O�����VST�xE�<���{mD&:�i�>&M7�f:��qd��έ�89@����K/-�����a֒׾��5�w�HH2(�M}�}�`B�fgg�c
�w
mv�p�=�� �%������8��22s-Lu�n��*D*�����'����Hs���E��q�Gq|��mv�Edy��򬩒q�3��?��ޠ��rܱ$i�i�x3��,���U��[�!�V�D蒫�⛺�B	����Lq`���ѩq*��k�Kƻ9�[��z�N�lb2��>�!��K�ɽ\�ޯ����<�9��a�Xk ��G�����8�jƨJF�Ҩq9"G;o��d��� b��c����!]�J�K/�u	'so����ҫ}���(���.��z�k���P!u�I�������ɇ=���p�BYI�`ۄ��qB�]%�Ex6�NX���r 8�b#&��<�������m�
��b�,�g-�*P�4������]G}�"{a����L��8:V��@�.u��R��y ��9z�j������h>�G߷o���6)8I�V�T���x��zח�a��3�g��'ðr�c-�lEVH���(p�>P�'�m��xn5Sܪ�v����Mc��M�}��}���X#Q'�K�D��Q*�����2g6v{��Q3�O�U��Z��-���aL�PB~Q��!�V��.����V�W���H@5iVM๪����c�u4���r��ړ<?�_���jx,%�����7(R�%:�E�I��ߕ.W//
	��W`��8�j� �r���Rg2�T���M�)1|1�]��>��Ӿ���{��%0�O��Va�����,(m�2��a�F�/IT�:2-�b_~��@�dv|/��"�4*���x!_��H�ɨc���Ln�PP��Q�����ѐ�8��v��߅3D��x����e�Ҍb08�:�JO��)��WL��W�9i��#�_��o �H+d�r�/�� �	����QJ��T�?.���ݜ:�
>������rH�pq�x�����.qC�e����/��+���7z��t)\#�t\��cS;��G��o�z���B�
M�,g��~2�#F _+�~LPĩ�����Q���
.���;/g*�Q�@8�k7���Y����VЯ����hj���r�ř��/� ?8/u�T[dC�{���dt>S�&^��{�:`uZ��	��%Ż.��W�8����>7�X���:�E��\JNBl�A�~�v��ӣR[_E�Qĩ~�lIb��g$d7�{��/�$��w���>kHv�?;ڤ�S��1�VR�V�9
:���@Ҷ�Xp D]� �Ʒ��Ht�6A�6���t?e�Cr���0bе��R:�>��v�!�R���|بgP���Id?ll�hw�^��G�,����o�]����]~AU�/��}�c����c�$Z�8u:^��}�T=�,5�:?���u�zao�a�1M��$_SdSPXn~�I{��íu]��g08������~���s��}�@P
��j�I�:(pΫy ɱ���z.f7ί�o�^d �kW ?���I�~	�C�ڂQ��S�q36��Jg2A��L�rHȟ	�=�'�ymgJ�BͶ�ol�5l�H��.p�v�[W冸��ob&2�<�p���+��'��ӼC�P�w�T��?�%�#Cv��c&���k���{�
�%�,[����Hs_A`���"�(��^ @����{�z�+Ih��*�w�EL�W��.�m&�wݩ��,������֊��t�0� �*ͽ��p�͕�i����[GR	5���K�H]z�hSA��ʦzR�͐#D��p��mJE$4FV3���F��L!�o��:�j��'���=3H"r�C{�{�g2Fi��XB
`��`�`�3Zz�lSG[u�ٸ���$�Lz;v����Й�>��-O��-Z��%��z�'�W!����V�Rm�}ʗ��'xzʮ"��\�Nw,�B_�t�5H�寁b{�u��\Ϧ �Ғ��y�ٮL�r����4af�t�kʨ/ԼO���Dݣs��͎"g��0'�!f�v���eD�h:V�l�(�@=D�cN�~�R�����I��wU��^��S�w3Xc�1�ę�0�=/յc�`|���0Cb�%Z�*��
A*%:��� #��	F���:�bdv�~;O�q��VwKw�����.��9q�;�9��ܛ���,
��/��i�p((����~���od��;q��O�r�pdc��2����9F��,�Q���+���]������E��A���<�KRجv���%т&#���/�nmi/��\;%�u"p��?��P5�JR ɤ;�Ժ8+eIZem\6�tmD7�O�\�ȪتߗBl��bksR� ���0�;�-�#N������3mi-}����q�iG�A���W|�<�isY����G������ �m<n=U�]	�#�lǂe��!b��hq
uq���Q+l��7�Q�ow	^�)�����Zv:UB���O����,�&3�$�-�Ty�q�-{��w�9Qx�tIQj���)"1z�A��d�D'ە�X_T0��Sm7��ջ�&�eW�5�
}�&$����dq+Wp���c�9UÏB�����F������duxA|9*j�=k����Ȣ!������'��a(�5%�R�o�e�8vn؎�H���q8���=aHC���tE ��s��XƋ���fї�ő�6�=?��;6yt���s	6ݪ�'��{���s�J��v�n�J�I�il��de福R����J6�X�B�9���z�D6��kd�~Y0��������3���b�6�X��<2��=TnS�y�z`b��=��r5�~k����1�ѵ�L{r�y��q0�ax�Y2��_���9�9xQ�G,��K�!�Ǒ6���T�%1�4�Up�f��q׹�T�ϯ��@9��z^�����v��Mί��ԑ搠�Gy��=��fm��T`�gd%N2с��텋H�"�u]�%+~�=��׮c���մ�����x��@v_{ �	K�=Z94��Ko4����e���:W�P9��/�X�k��Y�v�C`���P���hy�xG7@ ��a���}#z��a+�냒\�[��g�䚳 ��=��"|&�՗y[��t;ά�r�X}- 8/�!a���qs<Ӕ�bG�u�0iG�~-��%��̔{5��,�΀�\�R���Wh�2�O�{�۫M�O��1|����F�"�r$�k�G`����בmwm��hP`�:Δ����uK���eru#��5�>ؖ��_L��x��>Q1$o�5���P���;�ɮ=w�
C�A��6�U.����Att��u�@��"���f6I��los�/�(�C�1ȭN>�S���[S8I�(W~{�X�����Z�M�,<Ą˴�e��S�hǨ��h����e��*��
z<IA#^t��UDLH>�	�;�/ye�fܓ�}<�%�� ]��Ì6
�j霆Z����P����Q�4���6!�}
�|<Q ��l�c�+��\�*n�5޷�EDw��y<-�ņkA`y�������������H:	I�w�@2���.q�z	AKo�7�U��X���TBQT�b�*��ʬK9cyP�IZ�5��yOѿ"���4��/'kD���Ν�^�wt�'3��0�"����E�	2�a��eaqΨ������T�Ϩ��__ة������&�W�̧�Z ckh:�-�{K�$��-!�����
�5э�>�U�r3�A�q�F�|���ݳ�IX(׫�A]�4���:9��e�J��ÌE�ĭA��(�8]`Uxh!�g��ʋ�<[�{ t
I�}�M��1>Pe�殢�VX��?T]Su/!~ף������?�c D������j�=R�^!9v��V�j��N�'Ϸq�E\Cg�<*2��{0a��������=wE��Â�I�겗
1T��F( M��6��;K􋀘��L��%��q8�\>���뛮v�e-��Gs����C��G��)X��α����x 2-{�ni�\��	4�fb���L�%�g��7G>ӏ�V�� ��ՒL1Lg��\�Tb�U����%��D����=���c}�1jQ�Vj���:�SJ@Z�6_��Ƕ���亴���ï T���	�4�.z�4�ļ뱬�tZ��U�������{�Q�ie�ƶӉ)��N�=˟��R*�h ].���ĥ�U3��9���<�w/�	;�?�q2�1�c�9�/���'��D�t]��Pm����=
��+����'H@7�� b�� ��/�3+"d��Q��m��罪ƪ��i��g�0����Db0lو�$h��Z��I!��W'�>eqE������\��T��-)��V�oO�
@A��0)#C�,�}�[����|�oh�Xdpu��d8�9-���Q��Ʃ�n*�h�rH��Ќb�hMϠ�����#�8o�������({Wi��O���p/E�˨☇y��9AI+���pS��2�3�aK������T���� �.=}�e�#f(�\�����c��^/��Q?��z>�<�e��1��O��v
k��+��օ��g�C�F�eg۾"�C����B�GĞ<4���P��u�ڤ���y�.����?-�=�\A�]�������j��υ���)x?�#�����{���	�]��O���ɄEe{�ȁ����/ �`���@ֱ�(vkF�XE'Pʷ�;H.��l���'/KlxR.���M�{�k���E���?�)�[!u�5�(dfp��U �������X�ph�ґ�+�rpurp�?&K|2,��ukvk�>�2`�j�$�4,"�v
��?č��{��q]3�i�o�-J1{�9�3�PG.ꆞBN�	��h�ux��7�5Za���!.�Z�l�RFQϖpZ�+�Y��^���0d���0X>b'~F��=�AE��h41]A�j�`����8Y�T������m�ý��"���F�(�k�'ŘOhw�2�`���I��t��?o��oM�>9q��/zx�#���_x cN)=�x��f��z`r6���[���õ�s��O��D=5�U ���ّ����� �5&�r+K:��i����FwM�jl�!���F���/�?�x�u�V�T��m�ٙd�!/��6uO����an7AQ�y3��g��m�E���Mjq#Ҷ��z���г�)�����
A��f�N�8��{�����9Z��5�+�An��!���ۅ;�g��z�g�fL�čޱ�N:|K�i�ؿ����GT�*!�`3��Cb�������j^_�Ģ�(g��:=��1l�ɒ��+�?�����iXg�l-2x+�]���s���lh�&�&�i���1��.8�ˆ+ �_����R��!}�tܤA�x�k��Vg1g�����켊ovEV6c����5��kN�JN{6��H�ڌ����	/} !^�|2��(f8��5g�7ܹ�h��з��TO������a�N7�!�|U
�E�@<����mi(5tF&��"a)��vm"Hǧf#��H�6�����8�>m��������r�i�<�ü3.�����R��G҈������٨������	g�m=��C��f�J���@�OiJS7/`ᵌ��?�>��7��� w5���EzF�Zu�Ǭ�uҒ�#�;�y�w:tk�\"��π��ya���-����j=e��U��|Ȝ2&��f5�!�\�P�+a1Z��;$I���^YE�k��J��F^�&���������睱�#�3�̄�WN�|<�}�
�$=Rݵ�m�gOsh�._���=X��` ὇�}�$�d�O2m�#���aY�@<�L�<QP-0�t�wԎ����[揌�vx�\�D��!��c[�	�������>�,	&IDC����OݘML��P�'�W�|*e�F�ǫ1'���Zсl&VC��������}�i�[�}ً�@n>+c4����|���r�l~5����gpZQ���Ҽb.�-��H����OݸSL0���MY�l^�?����q�3KN��\�$+�"�e�������/�ޡok�>a���Q�&�E��A Ŷ���F!��tt!�Rd:kbU�Y�۝I����C�u8�q����'*/?Ɩ�٠u�n�.���\	��e�8R�ʰ`��a	��s�s+��$A�f��8��oKۘf�W(q;����Ix������qYQC`X����Y��aލ̆dy&�������O�D�b���|}�䶕�PU�����	��kJ���3�J����[� 9�|���v�`�+��KY�_�� �K�	#2��R�@m�?g*�nu���O�Z�Wx|�l7�t��=V�`E4gk���+�]=G�km�Z��	��ٗ1jp�C
�����M�	�&C�z���Jt�b(<���D~�R��W�|bՖ�&2;���� �i��|o\l�;�s�˺S�X[;�&���Y�]i!�cq�#> �vRr��Ƿ��3�5l�Qv���؉iU6��w8�&� �D��R����J�	(��V�l�� �2\"�>�� j��-q��;��WX�Z�,L���@τ��G|�}�It69��"���7���K���L+��-x
<�������/ۥٰӞ&q5(6Bt����ة]�ߖ�~WTa.|w�i���m��{a6�]��]�4E
u�����\��CMh,�¥�����e�ɔ��Y�S�4���¶�ʳ]u���n��@�\�cX[���rW��Z ���W��=,�
+�jM$�汯�X�O���j��%*�6�ʒ�����NFkt�Ts$ų��|�MR_k�"O�r�I,(E�
|�� �l^4p7�$���X���o��o�k�����b��[
��� 	�RQ)�ܦ�R+��K������E�����X_?�����~����y�s��%^����J`>����r��T	f]�8p��n��uY�4U�4Թ*�vu��ۯ�lIQ��ӛ<<��z���>,�$b�T��&�}����2R��Y6ޥ|V'VV"��3���d��.�}!%���g_7��N��fz�v��O�du`�W��d�O.�4"�(R4RxVi����� ���(9����*d@�(�)Q�M�ax�$ [΅�P�/�M���&����gv�0�6'C�+��S�Vs~د�\���#��H�����(0̱�������G~i�&��'$�h���Z ��/��7�H(��B�(���� ��2sP�Y�ti-om�g6�b�"b$��rǽ؟hk�&��0)���n�)��V�7V��HL�TR3�5��?a���]���*.j8�Jjpǂ,o�@<�D���]�8��(�k�%9Z��
]s�o\8~u�M�Y�O����0U��f��2W���]�cd�A�AV��@��K�VD۸��s���=�7VmeZ�?�:�唃�՞ϒ%����C9�y5s5?��˶�5�ȪB^�2���Y~�{�{/";d��1��M�B������Xq!�8IZ���>�7�i��a¼8=��ǎ@���~��ܨT�,aN�����GĚe9�$��P���;q�����U$��$�~XhT܏}_㵃ţ��v����JA(ꜴrGƂ���Ks^����唐Lϱ��L�����m�Ջ8H>c�̨R�Ǫk�bq��B�	K-���ǈ[��T��'wxٟ������J�8�e;��ni7%���L2�����ᑍ�C-��|W�O6de w���ݷC��@�Y�!�YU��b21����"�>�P@j{?c3�q�	B]ig
�����}�*c?���T��p�"
��u�������&)�9�7�Z�X���ZH�m4���uxMhsq��T�������9��C���%�U	=���K��2
�]e����NN�3�1�M�{����|Bԡ�X���'5_&g������kѪt5'Vqu�b����������8ں��I;08c��MȸD���/T{gILR�R���Des���ѶX;���c�;��j�W��R7�����x*ӬT=��˕�=q#��
:�����N����j����Í���qa��`riw2�p�o�ɗe;�D�K��p�>�u�sC��5Q[�|�,�6�1��:�N+	
��F8:�:�Ő{�E2��^	���|XiT=x+C�w�&�,�s_F�CZG6��s�x+����V���Y��-�xزzB����|�|;�BJ�3�a��m�?�N�B^��%�6A� ���
)#��;�%ت�{���x�	8@ѧ�t�<����]$����_�QqK^;�����<_}�0-�2��l1�Ψ^T��e랝a^zr>ۀ]���"�J�Kʌ)eE�h�^�[�� @���ڧ��(�[j�Ca�Բ�	��ž�FeL^Q�����┥dEN5�CUǼ!�mV�k1Y{ŵ�ǯ}��X�˾]dݏ�(�u�6j���GX���K����hw}'��ӬF��\}��������U$��[S��&5�޻��8�:Xɲ%gT�/�PV�sPu}�P�0p�
�1�@Ki�~ҭ8��V�����kí�ً0^ӈشA�5_�@i��\,~��2���K�a���i!pV�9�-գ[2�#��Cssf1����_D8��;�K�4~�]9��:��/�} k	�ƻpj%�%�X�7���aY'�[#�n7�٬�A�H���*rʚo��&�s�e����@�4$ dy�H|Uh�F������5��m;qӁ	"���'�T�;��AO�Z�;���
��~������"ҩ�W�	hb������L7���dPl����0�)o'���U>e�?�Ge9��p�	(���I���g%�ޭ#�����%��֧ۨ���!^�T�<#R'��cԓ"�)�/�:��~j�;+�z|�]�ݑ���yx�]Y:0=l�P&8�݈��`@��5-� #����h�pXŝ��%��I	W�'�1�n�>a������5sT	f͉�Q�7d�'BT��eXkeE>k�5R<Ցq��$qv�';��@��	v�R�$�+ǐdȞ�I���ڡ��v�ڗ����z�$I�}�u�H�Y��3�lq�-p�F�#PQgB�|�ؑ��v�r:n��R`�u-�'b/_�A̞P���z@��<2%��Gy�65e�7�e|H�kC�.���Y�mjwgU�6�]	|�_o����w5�-�0�@��F ��IE����5�����8d����՜eE�ޮ�0��%�����Ct��\cm���DZJ17�z5:��m)^�������v5��g6���3�/��9"*%�������`��[�Sz�+?�E�&]K�I}g ��E�>:��헝ae3P[Z8�I�i�ˮ����i�0��
쯗���!���݉i��DX Z�`�rm�(�ֽ�Ւ�n��$�d*z,+��6p��.O��|�D����^�����EE��8���� �H_�2_���[~�K�lE�v��l���L(H�s~����A�o��c6���J1�i��8���f��đ��)�]�Mw�}#������C�y�|���T�2r�>#�C�d��m_�?�}E��A9���{�4�
������]�L�:WX9��s�`�ץ^ew�����F���A�J|����'�I��"ȅ �Be�Ph�q�5����w\���⸹mL��l
W�x}WyzD�t�q��ƿF�z|O�!A@93���@�a��'�
�@cY��T�:b�t�:0 ��<�A���4���$����[=��0rhۡ@CF���ʝ��}{�~��az�M�Q��9<)�_����I�cR!�/��� Y��m���s�*��w�D�GC�笪+{=���Wļ�3�X��%2X V���T����;�L�E��3���
��zg�:U��o��<����T|b�����4sIYq�H5mZT:f�/k�&�S���#�Y�wkE���]
�U
��V�Q��^�e�L��Q����(VE����*��E����BĎ�41�T)�N���������y���=�"���/���vǏ��_.A+ai��3T�t��Q��RT��E�o\[�Lgw����:�4�ۍ\0�N�Z��$~PĈ�D�zc��~����������۬����-�l���7o\X�j2�����+Y��(�S�g�C� @:���[�'�g�_�6��k�Mr� �y��~뽿�0v`�'E�C���^Vtu��ؼ��sO��"��Zm�)WX��/A���Q�L�x�l�$�p���r]v�ѥ(�8d]�=� *[!A��'t��)���[�͗oM��>�Y��vP+n��j����K2��5n����dDc��2Q����YX�w���3B�'���oV��
:K���˹�5��s�+R�<S��0;�ٔ��\����ކ%�����o����%��z�BL��L� �IX�C2�묠��h�1ê�R.��e ��IZ=���=3�iU�>����o�l���C���b	!�O��;$ _����pՙ�4UZa��d��^)�}����0� �4�ɽ�rA#&� ���rY��)=ui�G�K��s)M�3�E S��p+p-�|�.�y�Kc�gR�ń9kU�iGU��:H��^�{tuۺ�@��%'5�M�0ϕ��Ր��C*g2�����Ȗ!A	2\�|���u��){���Q�ˏ�[8�#��;
����2�o��0Ѡ��9�2�[Q��D5s�
 P�NW%�ݞy?E��g�g�
<�X/���h�B��-���y�(���d擾�� k�R1���$C�(�d-��ï{)�t�aP��f��� p�����)cv�L8侩U��U
��}�f����x䐇������'�j�5�F�Sv���L��S�.�"a�D1��j��܋��$Ź{��.��7�qɌ�X�B~��na5��.�a_��=����W���t��Ҡ[W���$`6F1?0�/�@ڦF���YTE����ψۉ���t���ǀ��g�*��UhmB����%V����+����Tػ�|-��%�kH�)��\�8/��dÆGF-Q��v�G�h''���7�%׌���&Tu]��a���C���X�������6�Ę [����NXn]jde�V8rX9��n�q>�0�̒n%D֮�q3�ny���`�M@n��.���bYVx���K�o6�o�FI��E�mO-���,B{�Y�8
�}�˄�FX)��*���$	�U!�r�y�Vq�]YRT����&dݱ嗬��(����~�����u�Y������_R� I&�wJmkז+����㳝7aYh+�ĬHp��_5�b�{��y~�N��u���O<
 ���l���|��U���Nߍ��lP�@��b�@32�;=`��ӊ�ԭ�r?��j�lp:$����L�]롲/֛����!�2(�����z�#N���`|8+4���{�֒�x�'��/Pd�C��tj(P�ΕT�*�GES�����$6.�JKuI�P�!5(2�s��%��~��WRa��5:�����y�C*�k��υmM|�h٘���I��5��tT�!l��F��5j�-�d�%w;W��cw�z��C��fѨ���U�]q��@�.
\k�����\=�U��Zz,�d�?���D�w���m�7G�"�o8��=��4{��H��J(b����"����d�D��O�{~�����U�	Hm�#F8g�*g��.S�z+{��A����϶�'Ό���6�P	$�8�Msp�<�q�����v�+[Q;_���؜���.���*g\�y�O�1YC �ﾀ��	��\����ᆜ7_���C���� �Gs�X�#�y����em#���R�N0�6�O�r��|��|��?�
��^Z�w }\(����4�4�� 6K�1PQEAUD�`$x�U�K|"���q$���$���=
�`��҄�s�HL����־i��v���b��s�k�k됪�l�^|����~f�x�Z����ᖄ�mGf,4�T�21���PΔ�
���,~��|Q�B���_#�Or�/�I�r�����S��t����]�,9�q���&t����]Eғ�ݎ�^��Q[�L'ׄ�g݀�jH�P l�4����d�����,'R�L�ճ��H�0�H��V��u�Dá4�<��PoW���X��.5b���,�̣y�`���;OC�k�FȆw��p�t;+IݚNc>�{�?͓=9p����/�G�-�8p�:��zڈ�Y��W�ߤ���xwٱ�N��=L�4�-?O@y�|!5e��UYn�h�o��3�}��ע哴h䆙������g
�eP;��`��!/><y�<�:��L��G��������65�k!�d6��M�c���ڶ����^�(t
�����T��R��=��2��@9B�>fQ�u����ӟ��b�b.;+Z��9�s;��yQ�v��3[����*}��T�jJӄ�p	%�YP7;]�p�1�n`���y�k\�$t%����/R�Tb��I���1�l�&5�ȧMDbD��~7��U�:��1E�e�ļ�Y.^Ǥ+Nǀ����Ҳ��|��oy��#$�d���Y7�$�M{Q
!�7�-�(䉳�8� 8�������.�M!�闳<���	k��I�對	�d�{�5Ⱥ��H�f���"�_Qm��꘏r�{���I���2wa���e���5Nw��ܹu��7S{m��uHs�w(U<yݒ� y,�h��+R�B��/���*��9܊:���Y�L�2ٌ5�/�D"p:O�G#V�'m:��n*oே X�b���Z���q�"h�܅L1t�M�o��2�.0� v3Fv�P5]�%�%��⟂=���t�]�B�� a�o��(	%#h�Q+@9�4�n����Y�6a!�:�`�}&	�5���VfoC� �@�/�
O�����RYzd80{?Y��RQBR���E���?�����T��s�m��	sufq����*��i~��ЋC�`�ۀ�D�{E������Q5B]p�Ԣ��i�^��	G�^+��J_�;5�#��)�!(��(\�sa�k�e\�X��F�Sݎ���?��\�z���sz�e�6����Gv���k/+'��!l��1N,���P��GH���"�@��c��5�8n,��Eo��
Ω�y��V�,������w��w7�����g��E��2dq���Wк�<�.�D��z�	`p�bz�}�r�_d�ź�i�bĭ�+���� e� }$@�wX��Dⱕ=�3gZ]6�'�����U�Y�nb-�
��2J�;9����L�znpTșn��ѯ����[�RL�����x�؀�E��3��(2̀�}��9W��h����p�&aL�3����_
}wZ��c�U���Qv�x$����r^3d��1�-?V"P������S���9��p���b�4�V�K��ޡ�מС� �m�)�Y��v8�<��f������}�$��ou_�k?o�6M��L.d�C���PØ2x��MWL3d3�����s{�bnG"3#vJ]=�� Gy��z��coJ�C_�N?��[��0����PtE��q�)�HA�§|�䂅��eX�֤ ��6b���a�`�S�S�{��Q�^�B.[���8Z�v�""���E��n��=
�*lΔ%�e����c���֣��D��̕�F�4n��d��"�؋ל7q�R}(�������w4鉐� �)�Tݿ�,ͷ�E!?�R��S���`�U��E��1K%���H��
�*�s[G�5�����6�H˔>���R���%�)�v'�z�?�ݽ�h�S�9�I BS�pr:I��
ű� �ew�Ct��]�[�h�ч�w0���AM�>�i[����E�y������8�]:�
4�>�+9S��б��+ܡ���@B#���m�Φ��{����V��:����dT�-����{�"��v�l_G�_�ѩL�[�����{ћ�<"d���\�_�;��� �
������,RYq�0�7%�/��x-_�Y�J7�O"�ٟ�?��>��7�'V8�4}^�X��&�R���hm��2U>'gb֋Y��ۿ~6A���NZq�,e4�?����м�g	l�<܍X���F5�1�-v^a�dT�g��� ڽ�@I��k8_�HXز�F)Ad�Q廄�$��Vt�� �R.Ƞ���K(�sVɣ:�.I��4�j� ��Y:]����}J?�
ǗQ�����}f{�ojr�8A��7�����U��ůj����G*(����5%H+����v�6������	U�Døwכ��9�W�75�X}&�@�bbT��?�o�p�j�Eo7�0�\&(/$E���7����͓������ͣS)!�_����#qt�k$���Ǚ-ҭ��Ev��v��K���`�cQ����|��k{%;v�+���)y*?O;�g/JkW�@d�Y x~�T���F/Sp�^�JR=4�:��?���*��i�[��'�����@,��ޑ� |S�7~��h^
������'چl��W#<.nپ,JZ���O�|�S��mk�ff׫)�
�Hi��t�w$�(��$Zp	�E�(*�vaU�.��X��ʦ%�FI�KJN@a�[lPp��fd�4P���_�$�4�ȁ
V+ƂA��n�_R�ƛJd@����������ނ���W^I�����1�l���J׻s�@x�p!2dQ�	�Q����`�v�l��
��*&P S+~��Y��0D#�?�����O�kOĮ%��U��������ۨv b��AM�%Ww"����mzK:k-R����շP+�����~�m��Eg��f�ϲ��E�� ᳞A7�<=&�a�޴��k˅hS��$�8'a��5�nb	���A��Wu9*xl��F-J�6��[%�b�;�.\h����F�	U �}E���oW��6�18��ş��r�1�u��}U��qTA\�6��"������w�yl-k�� \���c8k@��JsP��d���A��ז(����f�Rm��{�+j{��D���ar��XU'ѕ�ܨ�c9���Y�쏡_M�JM�` j{��f����ۨ��MEpN���^)��tV���=�u���YHQ���� f�MH��61g��f�՚'���~Z@xp4�ۏ7K��+�2{!�a��ӌb���(	�%���o���-��&Lꮞ�����Zz�i0��펽\W�PC��ڞx�V�e�u��k8kNx�ү|����n�{P����{7��Q%)MWH3���ӿ2��7�e{*�CG���s�y�L�)!'�1��!�8����g3lp�~�ũ��m3(q&���&,����e�`�CCXK�9Qc7�9]������0M�Q0E���կ~�����K
�����兢����^��JW-e�%�n�$th�\���0��u����SJ9)�|�������e����*�|mt�������S�(�J�������Z�s��#f�A��+fu��3(��ruc���?� G��T��������uEJ������
cGq���*�k�CK�u�$j�.���+�Т�]O�Fq�<���H5,O��
�3O6�5M�Ga�Q����:����S|#�tr���f�%5)�(������"2 l�����tv�X��G�{����0t�0�6,V�p��2|��A81�䇰i
�@ƌ����qU�����Z\�FEfXw&���'���ǈ�D�!��9�s&VܦOK���c�.��}�s�����9#ϪUEa^����G�Ϲ�붥A��3�~���ڬ�%��6�;2�6oy����Y�u+?��כ��<��B�GcC���囻^���B��gMa3�_J��D�vA��Fm�lϐy�ߪ/�ѡ��c��g�Zԟ�c~4�Pl�>L�|����z�*�p� ��Pmo����>�1VE/c���ф�G��cm[~S+N����<e	JZ{�P6��MM��~r�4K���|Og1
Q��V��N������IU��O����z3]�e�k�Q5L +�۰��QM:|�Ǳ�?�l���t^Y�.Hy}4�=�%�,s�Q5&�}�R��|~�$L�@SWY�-����3��Y]s_.�L%H��K�<ּ{; O�a		��޷�:��Y���6�a`Ύ��,*Qw�5�1t�� *�����F�q��c�ܛo^i�K��!]�tq������� �kiͿ�*"Y�އ���^`g*�j��"��ky�E��h��m"7n�#�B>Axip݈�o/������.M� @lGn��g�s�i���*��]J�� ��_�Y��T�U=h����F�"F�b�-����p�E"���*�Np1�F@������$�n�3Y���6�h��d�so��l�`��X_f��at�v 
�ܓ��7	��v�{/�s�U��V��y����dFod��2i�T�9M��|(���tԡBF?IW�m���ˆ���9G,B!9v�V��3h�Ό�$'$����5�.(N�פ�t�@��û��g@9��&���փZ�Q*}�[�I�8�h�{+nv9xڶKO�F�_�P�;�|L�;}6]�A��y(��:|�������;U����L�[��<"��|��x6��ſ�c�أ�:����/:�i+ő�**�sWM���K88u���@��$�]W��b�|�I-ˀ�a������%�v A�l�����@�7�!,`#��/V�J|ճH��M���	n�,�B/��H+*�����",!��_�'�U�>��T�,�̆Wk��X���O^P��4� [yv��F�%:VgP	�w� 1�M����>�C$M���r�|.x+�K7U�U���hQ�~_S�I�XxC.E��s����2ԫ�?Y�[x�S��ic��.hDz�:�T%I��rd��O?��P���c��1��1|m�-3��mY�n�Ϥ�~���:����5��
I$kN��#(&8.�0�w>�H�H⻫�%&���K�����8���a��=��r��׉�Z`���_��NX��5~�6��8�n,�v{Wu��d���UЅٓ1^L3�R4����rj����#�W||�:'�m��;o*�\��u�=��KS�n}��	��G)2J����K�r��#!d��!yD��@>a���M'��$s� ~#�8�L�� "'T�蜌�=�dw�+r���&a�7#2߯�dA�~gz�,o[��Hʷpch~e�	Q�۵y(�Z��x��8*˻��N;
�5˩(��<b�:K*!��%��Js�3}$�;��&Jκ��/Q�,)�"�q��^�S3:Mw9#���~4��|�K�L�W�f���vвqE\/�`1B_+E��9�ĕ����lN�5k��B�$b����|j���RT���!��K��0�6��P����{S���I�]= �D��	+/,Ƶ��E�g���L��+��. �&	��^y�_�]ײ�GI��\�~wy�#Ʌ����#{��J����QdgIz��ɣ�~�w���j�ϳ�4=:ZE�6�{#�Kj������)�&�ּ�==�og�oƜ��	̉�r���B��>��O�4��^C`Xh	���2�IL:��AAM.[�#7�69%V5�6�ݑ�e��Z�SC���%�RJP��`��؃����������doߖHߘ@�࣭"A\/}�.�u�Qq�U�	�y�1��A�:/����D�h;��$âe�)�kh��\x��H�����6ra����'h���rD\�y����T��������a��7�ѻ�L�����\�"�]�0+����1O2x>f$F��:�0f7O�P�����	E�Ԝp!�\�$o[��}��"����#�����d��ۦY	B.F���A	bR�W�x���O���q��a�߮&��]�����޿Pi��bG�`9��+��'c�c��'8IS�ҏc�ʫ�O��?��V�'S���ES�}����� �G|�
��YϾ�����G�5��T\�O~�tQ����#3nSj2�0�j��Q*b��#���H�|5OM��F�`�>�)eP���`�s�&r?[N��YfvQD՝J.qH�*�-�W�x
7�&��җ��J͵���ѹ:�4F�{��yQ5�gI���h6� !5B�m(Q`�¹���k�O�N3!����^�#�%k�KOF	DP�+�6:�95��	�2�Uɂ���u�q*�?hY*.��{�0R���~Q)��v$f�'��j��#��DS���s�@�92����-.�3��h�a��ot��n'���޼���v�?�p-�I����f��s�2A�B��Z{ož$���QU$H_�~�����$E�
q+S��ഥ6H�P�d��I�ͱRJ���x��o=ShO|�:�`;껅0�D�I����q/�/0�������� �CV
�KTk2���b?�]�A�+�]�HS�k�C�/"��Ht2`QL��5:S�n*)whzϊJm@��f���3A��Ƌ-�h�;�S��7wIT�d�0&�Pm�e^6.��Z�&J����c(92�� �Gb=j�ղ�Ŵ8�<Z�Z��k�v���.E�f2�Y�bI�U��TAX0�C_��k����/�].w&K��]�qɅJQb�Qݮw�}@+��R��U��%�����Ocb�rG:$�Z��z��*�#��w.� ��믵Z� �B=1s?{2]��|�|�!<�t�eJ�A��1^e�RA�����&��>��������+��Z�_�-�y��]���j�B�0�@�8��#�-2VD��s�:�F�Xa�]L��?�����^���y�)2��w��ޒP�L����W3���N�Y�]7��/%�;�`�6IU�C�>�w����J���?��IAȩ1�o�c��iI��I�^� 
1��q�a	����D4.��T_ވP�,dY\+�ӆ�^�'Pw����&������ܐf�E�F�k#��&B�������b5ǫ����y�Ej���x��O`�#Jݓ<�nS��b��1I�;YL�BM��{̒|.�$jU���b�����h��{�3��� ��L�8F���!�KY�iG	d��d6��\Aٳ�q�p�*/����.����؃�_@?�Eס���a7+H���m��`@� ��Ys����w��LUc�$��WђU�(�I����$���z�)��cR��[k��TY�^����E�D+3�Ly��s�V���A�Þ	�8���3y.ORõ�N@���/������Q���
)yߩA��.�s�������0̀+�������s��I�q�nuL(��C{v5.c���K�U�'����%�`�l���HN>/�Tf�r,Ak��l�$�5K��>�a����ۗ9h�;�W5DT|P2��ϓ��������!<S�עٍ,k�d�Fd�b~����޶sWj��ʣJC�����_�e�"ϝ��i�4ζ�#zYh��u�j�����a�������R���<s��H0��T�ɏPY�>jB$jTA�(������5���$��LF��-|�T>�7�{��:�ٞ�x#��tɽ��I��d�s��T�˳�~UJ1��k9ჹG ˲)R���^����h�^�O�����Y�����N}^�پ���xg5��I�s�a��p��|��������o��D��	��&��5�6�II!�n��h��jߤ�"�$Pּ�;,��qF�BK���x(�~���v����<H"�8��7���|��l��2~��q���\�����N���XP���9�JctƵq�)=�:ڋ�>���)
&��1����L�	����,��/j�"FЫ2)}F��8�hn�f����:K��:�i��x�jU R�+�F��i�� ����~��ʻC�J��v�#����ʇ�.��)X�ub�pk32�����<*���Afo�Km�oa)�H��:�|���)����b{qC�b��sa����,d��l��UM(F7����/D��(���a���xx�Ӗv�mq���K�y4�3>VD�pTR�kg�H��� �on/�~.K��,��&�z��D�GQR��;��Ӵ�����,�ޫ-�p�ė�l�x�)W��̪C�H3sN�Gf��	Urh䱁˻��mw�ɯ�u�_��Vn�YM"[��a��nN�{��gZ����}����P�w���Jb�՘�p�MCѫUs-X9P'e	"W��@ �P�\Ό�ڵu1Z�`����E+2M(�'p/��e�a�s�3N���G�Z�E�����,�g8�;�5c�2��Z����ģ/J_��C�T��lD
g�S���6<���˗C�M�7[p��o��L����k��Pd�RfcC|1��f��Y����A�1�L̐LKVM#ԛ�]̨&"�ۘ�,�3%�<hı�#�~�Cp9���_��85��%+P�-3��B$ł����:��Ř�e�K�
L��X~���u&ƣ���D���
(�3;��7�1�/H���Ǉb�P��@QK=[�7k{�?e ��r�?���3���	Z��H��w��K_�x:S}��h�h�e��)�D�y�:A�3����<�n�`�[�0��'�v(z�LҮ_I�D�8V�'Ӕ�)������	(x@/G�E|��/�e���_��h(ؐ/o����ӗ>� ��7��B����ģ�����d��Zp���/^�@ΥC�R����򬢢�;l�j��Q��B;�)?�Pj�QZd�s�cV3���R^�s��Ë�,��>�t�)���Z�*�:�n�Ԟ���MXWQ;�\,#x\��O�˂�h��J�����7m�Epf��Y����>ս�P�
4)�j�d;ĉ��Cw���g�~�⍢�5Q�p͑J��̂�|0-Bz�����Fjk9�{_c|�w�Rz��	Rۥ�Q�x�t݁��|�Ss�����9�g,�:h;�W=���Gչ(j�����ґo7L��	x�3����u����m{�j:�U��C����\��S�x8B��e{��s�u������������z��8� �q ���&�0�]FW��E�A;�@����0۫��3��O�Z�-��(��z�|��2s��L���f�V�k=�����P��-��լW��=�����"���5�x�����F���B�����!��IR(2�m?�S@0��_ض��u�U�@
������[�ڏ�K�)Tsʗ@�̪уJ��58�"z� 1��ă92��ҏ9y��gY��.��3�)���Ί���iEz�<9�X�2��{��G]l��]�G���i��,l&��I�4����\�?�7s(���L�.�c7��}lC�o�{Nh�鬗�)}��z��%�Lvi �E��n���a8��I[Uj��~���'�@q긳 7=ⱝ���z��ϧ,Ȩ�,������I֢x��|����fx���M��;�;$xVɇ.n)ӖG����S=wNl �\�h�~VK�I"�M(�H�7C������ռu8c��w?�y'�'J�!�#S(��c�"�6�{���]�#�����*��FT9��FP�s�O��m�Fz��`��6=��@���W�8��M���b,���dO�d�J��x���|��'�D��j�O۷ j{I+e�M>M��f���� y0	M#��x�>'e�����̳�+�21Z~)C��ÿSmx."̪	S��ձ�1�PV�0ci���;�݅�;�)cr"��[d�
�]�X�Bz�cFa��� ��Z~���8��a݅�Y�n-yV�g�$~�-1jh�KP>M�A�dF�)-w�`���ѳ��c,$p{@�*�� �R�����U���<��tQL��	��d�HV��e]�L � ���y�����n�4H�{�n�'��m�e�䣴�x����N�k�`cA./���}��oˇt��vB�W�>��A��j6�ObA�6��>�s�L�~����X��|`�O��b�,�e���p�K�gѡ�s?dJ��m��ӡگ�o��F;/v>J���v))%jKT�.B1�!z��0��f{��k���e**{��C�.0�˔�G�B��o߰�X��;~�p�L�G4.�,�#���q	�����5���O�xs�ĕ����:�z~�ekƊ"��x�`w��Ieq 5|�4�z�2��j�q���%�i�o^l��4��Zu¸��O�&�ݳ-�}7Kb�e� ���q����:��O�6��R�Y��8�/�;�$��_�xA��XPG��n?0�3n/m!�������5���t�����Uj�����%�Z�n6�ȶKǢ�s�M%͙Ϊ���{ת���]��<�X ��TbO?��g;�H��Z��u�)h�?��ݒ�ċ� "�%%��@��ӛt�Ũ�z�d��jkN���/o��D�x�Qp����#'{�'f�.���J&��Z���2@
�)�O��(�Vz�
a�Tv^-��G1��^>EE�e���@͹����CGw|�YJ]-Y�lu:3(�
��͗Їwwh;��"`nE�ڡ�n|:I �UK���D�R�0R3���N'A�K�����Z�g*=f�H<�ڐ�g��f׉��}f��;���+]�+聺UE��r�l��rU-o�G�����������-ˬ���F[2&:�;�^]������(�F���Z��~�k^���8��J��W͘�@�����w$��QG���R���Z�R1xYq�=sE�D�����������;g6u���<H�h"�ƶu^㏂� Ha"y�}i�`3~p׊�ZϦ��_���z:��`ғ�f����Eύ���}��Mn�� |D\�8 �n��<��o���3�����N��[}�9x`x�"�g_}qUB ؉�I��`kR�]Y�|�,�&�O���ӏF��1}���7�=��ą��Wx�69Ot'c�f)��3�Pwa8o�5Y�B�+�
KE�pഀ׹h���L	��߬1��ʄ^�m�q��X�E�n�P�T�����v��ld���-�{<]�14*}hq�Z��*<�)~񉊹��1�PZ7ո�ἡ�x(�i��ę,N�Dݑ{���!�\��6����-dU���I���ij9�X���k9����<�U��Wh�a&h�Ӊ�8U�5��4���8�n�"��<��K��~]���H�U�Ȟ�xwg�)&����h��t\^�ؔd �5�Վ�JU7���|Y�ݿߘ��պ~��W:�~�"B)����:4Ӛ;�;��C��X�w����˔(%U!J�3|��v���$�����������|��V��L&�bo���+$����+�7��M9$�@,�	��T��ڪվ6ݻ�Z���v��d�7	��$	ʗB=�G��	��z3Q@���X ���=�����>��WU�˙1��wՠ�B��ƺ�&�]��+�ݾg�	�8�>߅�����7�ƥ�/�kE��	B
�8�8~�/�^�v�X�N��#�����Bл�;47���<��:S����=�~?���0�N� ��)�d�#����Y�lP��A�}�4�n>l�rxLd���F)y�B�6���a�L��<_;P��H��d n��0+x�Y!&Xs>|8���E��=d��A��X��d	����0@ZU&;O�r�	�!�;�����29�z�ȑ�@���ԏ���x�K�T���L��^�me��`���J1{_:Pz�|�W���o%$G�.��Y5�ܿ��`#�ߵE�Ӹ-HF�П��}Rj�㩘*��H�SnlORvu�-��m�T". kۘE�
�+���l�����s$.d���>�������Ӭ��L[��@%�J4=�Em��S&՗0�����１��S��J87lƟ��ί�M����w�̛|���~Z_B�_�y������i�J���h�A���J���D���Mg�4g��1��)���:����!�]DK���#]���Ly��hl����$?��wN��/��=J�j�!r�p��M4K�U�C��'�=��X*�:��R|"��69�	W���%�W���)�	��
^+�G)�����f������p��_d��6F��p��i�����@!e��V���&���2@��E_�,�p���"c�B&t	A��n��� ��Z�ix�QWqI��ڜ#߀l�8�ˎ������������a��?�|�Y �����.�!�Q���9{��x�����K�P|R@X&Fŷ�\�E����oT���`#���-VD�[!?��[)@7�m�m�����.Q5�~\_�t�x���
�zˁ� ��J%�t= �4یp�������mτcr,�񈍦H�������H�[�nc�f�~�<��07�?���M���6���d��EEͯR�������b��"�Ѭ�q��,D؉��"Z�I@�>Bg:�����0��eB0�ٍɢ
�ж�7����}~b�.I	(�`⼋��w3c ��s�V%|�5���������4+��y��c"`���n�h�)�����PQ)�mis&�4sU%���(U��
]�(�n}d��@�Қ��sj�C�L��U��R��u$T�(�v.f��@��=dw/�Az�3��FR��.� �FE)>[��]q�4�� }�S�����DδR�~�a�:���,�mf(�0��
a������U�<F��nT�x���C��(�E�Ps�����{�cz�����ogE]��dy����8�;���\Ma�: ���n7n��g�k�G��o���IH��Z��H-��E��e���ҭ��JO���H��SU�βWh�j�r�|q����EÈ��!�}*�-D(��s�jWW(���<�߀�a2�L�V뉑܆�+�Hs˚��_�mr�IcP!Y�2�-m,��9���>��ҿ�R>4�I#�.��n?�_;*Um5�7%9����N����C0�'�%?�2b܉���N��\>�s&u�\�e�L��F'�T!Sh8�������d���h�o��we�4в1t�"c��w�%�w�Me��2+�o\ȕ��+C���k���f�@���vC��!�^���_&�2b��,Z���R�k"s��}�b�
{�񘬦�����=[U���
Qe%(t���zq�;�����oR3<r)��h崑�Ru���3C4�xI�:��8t�tba��Dw�р<�L��� 3����٪$��r��6i�6�\�|�<�\��|�ȸ���<��;�V��i�Pk�ݙ��FnpI�.d�4�N	��rL�AOl̊ۼ�1��,g��5aM��(d�2l�$qC4M�S��y��9 �K�Z#��>�.WY[ʒ���IB�� �%��y�� �}�0���ʆc��P�^
�q륓_P�5�@裣�x�ɋ��!�`Z��JiSS[Q�Fݖtr�V���a:�۶3~tmCpd~�1�	`|�L�����6�t!�_Ǵ���~P�W�ądYn�����|S!Q�F6v7Y�z���D/9䐾�����Y?:+Zտ���#mrP!K,I�0'DAe!Q��QPyU�F���P��q-R����L�h7%-Z�`S��ic����̰����8x i0i��K�����U�+�#������f>lK�$1���w�z�q�?�w�)��/����*��*
�4L�.��g�
�|��ַ 9�t�-�%1��9?)6ΰ�F��SD�<�UD�w.l�]=���^�;���]c�C�{)��(h�e$�.�R�D�����r�1��͹�����i2�z> e���Ԛ�>�bTw����r^�E�j����-�iU���A3b4F�?@��lk{)aqvx�ν6�g�hV�k����GLmNB��~���p\ڔ�O��*�0{TP9�B�g�͞���-��+�ӂ
� .�_=��qi��ޚ7�^��-�:U�G{�����v���r�@�w����w9��Z"�O�S;A���٥8�X�$_}�2�.��*O��y^
N_(k,��Cqzkk�텸�9���\xuz���6A>�`�hIX��嵴��~��Ä1ϟ	u�&�j�!}(m[�P�L�����U`��zFv�qʏF�'�S��{Q@��K�&��t��BS|?��[])�W��	��e���z7n�Tt�2�v��@s�� �}B�����5*��2/����8z���p��S�O���<�P��;E[���h�a�O�I|�����w��4��x����
��
ke��w�<B/�{�X��\GET=�I#�^)�I,s\�p���G�x�nC^3P��~���Bw�*�-�*O�e-���S-�L3�!JZ���&�)Kck,n&��mڌ*�����p����|�����RS:�W���S""��'�w�ڽ���s�Q��Gm=>^���>�,g��-.�6d�`>����A�Eu��+�)����J��x^��J�+kR�U��Y6�nB����-��9ɟ��`�xp���\\.��-�����ؠ�1�*ZUs"����.�;�nCl��1�y1Tr�%F���h��ǵ��?��'���\��Mho��e��1�����NFU�[�D�Lr���C*m�(�,;��l���zB=����Ư��=|,��S$=��޲	�0ج�$�^js9�z��7�9kp�A��}�:$N':#M�A����sw4Ur�ZV��'�����+�����ƠX���:wO��:�Oz�����4��['$�FH�W��O.~�����d޸US��_r��B�S�qrc�:o�7
�R�VQ*��&H/ؒ��cW���H7�2�սA��g	x��5r�����Z�)��|��Ѕ���+��-�"�����X��?I�3�S��E_#*�a����l!-):GC`�2o�F�0��i���|���1]�4�sz�$lK�4�=3_�utU:��V���%��&%�VS�&�pA�D���t�����0��>�	�+�VU��fa�h�����&�H��4p��i�8hc��I���k�h�C�R�[�.i�����>v�bo�XI�r��Y=��G2��?fz�2%���� 6����7�Z@�D-@��R���*8ˢf�ݵ�!� 2%t�g���������x,Iz��7���M�����7p�L)#}��h��giH�]��0*��������`0j�G��<�����ӹ��h�q���ψrl�AT��t9��a�{2ʁj]����"~�8Jğ�2G���j�����f,`��_BŶ�R��H�C�ê���j��R�n�P�B��ޡ�?z	�A5�QHUw>*��R<���-���������="Zg��+�[�o����Ѳ�L�@9����&��4�8��>w�WA	��|J����7M�~�?h�����Ρ�ܹ��\�1hG46���dп��n��N�R\�)<����%����⪠U���H)��!�����C|�X�u�����GK��AO΀�h�� 9LWI��T�Y�;(��6�w`~������^�1�.���I0vU���;S>�m�0Ď][�ڲ���%a�;���ZF'@<ŉ�p'�x.�;Y���,�h������XM��t��"f߯��|,-�pp���*�%Y���[=�#��OYX�;�Ή�i��W��↪	o�~���[l���|0VH���R�!)Y�z���Eza��.�ı�< �U�?�OM�]2l��j�ZkJ-���������HW�}�?W`<.�噫��.�5� ����I�o [��_�w�`��C�Z̪t�A���oG*.��.qc�|�O�*W���%#��(��	�U%�Ќ�P�����D6�4\�h��ax�.wU��Sp+��p�����p�? �����Yl g��ɌQ���f宣py����6��8��Y�
���ʲg�@���@������vr�Li��,}Ȼh-�Ѿ�<���ͧ'9O"��~_j�W���eqZb��c��B�\t �Y��B��1]�����#�ř�e�� 2�3{��)�8i���+B "�<��N{���'T�qS����Ұ��
�7&�5i���n��
'��q��ʌ��ǈ�*��G�lEF4���$t�{�L&���������Q7�HT�m�ceCv�"�k��Q�:J���$#�d��:|{d#[wے��>�����܆;�	E��˓F�i��.��J�j��=#I���k|�6/0=��.��B����+ċZ[,�C�����SLk#")�A�H�bUѳf+ʓR�$�~��]F�0������}��wc�R�w�����\~$��be�Wӽ#Bxn��wz�u���uƇ��xi�.�V����������+�ƀ�����D�5ԀJ��?�-�}��� �3;]0�x��n��ܾ���'�QtU�1$�v���j����r��d����,�)��UOS�k�4�0�40R�Sм��{(sס'Y���K�&�l<07��*t ~�
�Qs��F�qг�\���VK�Ģ��T+� &K[gXS����[�ɖe_>+J)L�:�/.���D��W�֭�ƾ,râT)R_�cq��BBt��_n�b��_+J��v�|H�y�'	�G0ʄt������w����W]��]
&����&B�n�]4Z�m�8iwu�P��:z3F�/��ކ�0V׆�z1�8�3�� ��ioş>H&�<�,��Uѣ�fe��ʀDl��M�#�[���a�8�}�E��74��%H����MZ-�뺈�kcK��aq�yBoSN<>�*~lŔm��BF/Z�!�~�=hX��ss5�I�S�sS����W)���$��:ܢL#���-.st�v�pd��NZ�<��K~8J��X�/�_����?�dk������P���
� '�P�`Hh� ~�nP�;�D�/�,fn7ga���w�}B�=�I���� 㳓c����YĻ��;"���;XK�cL�*pHD8�, H��s��1��JA�0��?�����m�)�D�~h������\^N�xܧ� ZJq�G�����%�W��銮�2GW�r�a��2�YO��W^ð�O�Z@����6���&�9>����ne3"h~��B�#@�FKD�;�rըX��徕����9=����Z�#:E=CR�s�pl���mZX]��%V���$�dx>��}U�?�c�'���f����m=r4�o3��%�`��֯(������XN���x�LQ�h�Ƕ;^����������n��.W/��q��$��0��B"�iI���hVl��ƞ�>���ֳ��hw�F����!�)����s
I�[�r�s9A��P�s����s�@,�f'O�����[4e<���]-� +�">ܒ�+�MhG�>,۾4ʪ�=,Zk{R�&Og��=TS����5��.�/�3�c�H���;;9��ך�u��"ޥ�a�wK�rlF	�7�uik��a�ϵ�{d�(�#�u54�TX2�M4��.p ���̵���fM:��C;{��^�?b����i\��NT��z;{Wa�]t/w�>+��9�B2��ҧ,A$c�����.K�^��<�t��+XoW�>!Y�We��LZ-g$���!H����H�̈����Ɗ�һ0�'�C�Q�G��	���'�AەP��k��vGBb�
�7������rc�ꧣN�f�(,}.�< A�����}I�4>]�/�>a{V��\�ř���3	9]yѡ�=Z�1����m���pI�o�i,��mzV��ڔn��ˁ�w���x	Td"y��7B��z��]�{�1LI��k����a%��̋8��~X -�8�/h���{s��_��AY|�A�� �� ����t�c(6'��f\�Q	䁵rW��Y�ht'|u��A�ݏS�����!�6Ο3���>Ǭ���X*� �u�e�͢j���`��q��$���Z�孙:ow�l�t7�c��	�+#[�쩌�גH0i�d��U#��{LT��k��
��d��K�u ����{΁(;�a��6��� <�Z�U?��7��³6�H����.�Y��4a�1s�b�!�+�C�>�?"�u�Ag�	?wCwнA�ƤtɝH4�;��	�w_���ѕrD^�5�tE`@j�����vW���'h�{�{R!�W���`i�K��z��ҡj U�E�������F�N�g�x|-��va��Ɲ	�tX�T��B��ݒ��3�&�ItL)")4�@�GJE��PZ�%�h�<*��#V����و/���{@��8f�.���I�n�3����J]�������Ⴕh��&�Â~�H8��v���NN*��ۍ7Ϟ@�9���N���K�����dr�p�-y� ��C���,8+�}��M�nE������������n�6�e,.�W1P��|���}]2;,L�R���%}^Ny���"�bAA[��0%�F�r�%}��(��q���\��ar��.��7eͿO��o/�Y �jTa��ן�P`���v�e�V���B<S/W�z������d��WC>F���f�tP��M�5Z�m���'?�R3m�) yp�bqׯ��!���,J�uS��Y�hP���ډ�y��rUѺ󥄬���1&ǻ�S����Y���7U~~aE��ƶ��
e�oI����a ��A
N������f��mܤ!�1s��2�o*\k�P��8C(�A����(��p�?@��� ���{���e6Bs��?:VD�F�`~�#�u!B&4s\U��>ɛ�Jߒa@�8ň����a����X�=�2�;� -�<����;�t��8�`Ig彼a�X�	T�H$��{����U��	��=��@d�}���0-�'H��bjbem���R�΢0��V�#s]ha�^2�_�1�~��S����a�V�c�;�ׅ\�~e�1& ���Z�н�fב8ACcX��xT�ߙZ����;Mj�>�J�p�Ѷ���ۜ��~U�bM|[�}��K[2�^!�x�"M�"��ω+�\��ٜ�����$�ά3�7,u��\zӼZjEU�����n;�Q�{6Q7�XQuK��T)U�:U��E�o�p�Md�Z��ݑ*��2���s�m6�{AV�\ʲ�̬�禔x�(T����]�9r�����1������4�vf�2�%��l�\�]�N��.�� L����jO�T��#�����0�����/�\�IIy�,$}��r0qv+�mz��! �j�ys��;�<���9����j�Q�� ���Y��
���J)���t��o:n��)���{�ᤤ��ض��`�f�F;���� X�X2d}w:�m����t6�1�.�87��4��,��f$ҥ뼅�,+�[�W;l����Z�]Y�lT������(�KcVh1JQ��:�bN�n\��t0]\g` f��k�K�z>m��p)S�(R�������:�N-��B���Ǉ<��*el��H4�$K�\�y���K����g�GrؖgG_G�WVVQ�����] �f0�(�q��GG�ë�DU�)��qy�5	��"by	�tY��c<x�+SZs�K��� �d�z�q����I�����9y�%��2hfh=��(|t�h��B�V5k(�;a�g��Ǘ�h�z���S������ fżť��Ul����HJC�513}"	�\f��ħT�;��_N���0C�m�P_��b��U�G"y�Ь���%*E-�������Io%<�Ɵ�-~U'�8���D5}(�|�'�E���a�"i�n��^�=d�?�wg;w&��=��N�}������P��������\{p$�llS>���.�v�.S��O�uy;���Y1E"7���+�i����(��a����c o�ĉ1��htG9<�$�2{��dt���NsN'=P�.W��p� Gy(|UH���*��ԩ��.����vy��3�}J�M�qԔ��ޠ�{����`d �e�`rGh����7�~�����,6Eu{3��5,"D�op:������o�[��D���$�dc��P�a�0�gMv�x�l6�
9b������b��������6��*�0lt��j���݊� 4��ӕ6�ōd��a�٦,t[Y��:3���q�Օ
��:�*���(������9�S��g�o�����E�?[/yJ'�O1��yA�#|���J�	rå�l��[%��jȃ>���&��F�((���X����dQ��W�dp����.�,5�S�'1 ��+��5�g�w���n�Gg>�����Y{�NW�~��O��SW�LI>-	���㵽v��!��'~�%#nd�5*�ru-
�UM�=�Wi]B;�=o�J�T��E�Y�-&:,4�Y�I)���	Bü|��H�l�d��5���u������R�=������I�4����ˌB�����2�I��OB��b&�3���6�K�����OhV��b0�+��z��qhΤp\��+�x�%*�KӐ�j�j�~+�UA����8��ւ�'C�Y/1+]#���VH�n��}�O�Kʩ�?�R�My/�b�Gb�#�%<f���	��m�i?�V�Է��q��gu��-���	����1g�C,k�:��x���tw&b=�]���2����P���lګ-��]��O�:��Hi�y3�#��rd��Z1w��c1�Y�h�F�N>�PӾyG"�O6����U��{��	����S҆��7����n ���'v��(^��+����%���ۦ��mO�p�stu��>�(��� �*�!H��'8m�����R����@�_����Ԣqˌ�C�����H�����z>%YC=.ܭDG�5A�Լny�s��r����[�^Q�1�����q�ؙ�o�l�	�cUD'i\.9�t������G���P`	�t=Z�<��-*L<
<5���ɮ�֐���/�� ؽ�g�j.�sj�"��>�a�yUs�?�8̟>�#�gXh�K�gn	qj�����m�w�)G�ff$O�����ڝX�l�z��_�?��pŊ������~��G`�@o(�F��6cx��S0�4�
�jmM����o8f6��.�
�ϫ(��6vA7�9�ɻ�'���Q�wyf����E��}�'���pz��;��;펉������ ��b'�J�4{�dpFpˊ�����]��)uQ�uΰB��`5?��8G�IQ�Q�v6e.��B��o�0	�DTvl#8߄��1��gM���9�]�p��ݲ].�˔ƘЩ�A���,$e�#f��^MR[Q�kH���x7�]{�V%�~�# #�Bo[\;��p湐�[�~���K�*r;�a#�g���D:���X�B��:�)[\����B�*p�j⦣�d�F	r�,������mn��c�	e�@��9?֩n��B�>(�PV� ��_�wѯ��=��1�w����P��j��|�OH�wD���a��+D��:��K��4�B�׶K"�8N�h�@��^�J���C�(���b�F�@�3�Z�gM1�z�ĭ@d.����W��6?Y�4�Y��/i?��ܽ�>�T�
�GYPt*C�%g�ENb+���!TE#*w��+9Y.�w������T�~9~<l��F�$������>(ڴ	[G���>gٍիo����=IJ8J̼��v��ś8��C�x�*����+�EJ�֋��{��7~�h���O�	�{������@&p��ve��3�$�l 2��_6�W�;�hƧ��#��N*�(8|�$��ޏ�Ez�S;�#OÀW"��p�
˜ NY���� 통Tg�ǩB�<�%9P�UB�EH��%em���z�X_=Y=Udh�ӷz�0�C�aǥ�R����<�y���Y�T7�����1��b��
�:"ڑ�%�h���C�Fs��a|+9:��߃7�!�e�y'��$���!?�b��uP6�I��E�s�^
w�e�<Io9�<˭��A���"�xF{�6�A'v5G8�wӐ��{��I�A�u��EQ�P!QP�|�R�J5���ޔxF'�y��4X�����m�:eD�Ȗ�\��cq̢H)1{%	\�/-{]w��o�E���uk��9�o��N�[v�aT�6E�:��9�-�:2s4jƯ09<=D�y���'XL�J	S�g���	M�f�o8�&{�=������ւD�&�R��I��_�t�:J�=��#�U�����O�T�g����۱�y�҈W#b\��+��@�i���|��ɣ�w ;&�����Gp��[n�HN_�ͺ�3_��۞�4�ך㡓�[�V�����	�	����M3E��?x�|߇���6�'MM.�r/ �������@37��vr`�x=�;�n¦5��[S�Ն�݁j5a����(M���~�ϸ��M�$HX�$E���Y�U���Tƅz�����h<:	,W��J;B�[�@��kjN$9��"u�5��F����$  ݲ7���}�W���K(dKd�աb�t���6ӧ�T�{��(�h�?D� ����H:���r�|��2QP�)�𻍦!�Ы����͌=pRg2�҄��K+Cf��E0�8UZkͥڟɴ��0F���e�1��xz�z;N�uѡ�G���O�����@"��$d(�U�5����z��y tք����7��fL�r�t�i.��*����ep�#�/�RV��_]3�X"_�l��/�XE���S���p�)��6��:��A��6��'Ԑ>��N��u��Y��$C}`.zy�52�q�B|e=���kc��&�&�_J	����s�|#O�#		fuMeA����� �7$M,J��8�~���oo4Zҟ|)�lWK��ڮ�DN�7� �>=�����cB�u���1�\�6 --W�n |e'�/ �3���ڷ����'��K�<�B�}<�ݫ�Y��k|j����&���t����y5�w���L�t�x���S�}|6.ѱבa�3����@����Ƈ÷'K���Yq5�7QF�^/1��9+-Y�
�D�NԬ.��O(86A�LN-O��E�Ա�ڣÎ�`�9���P���k`�Jd��{R����#�If�xt��&���~���pשFEV< ���Fb�v��e˝��=�>���q�=7e�w����$�e3g��a�U���<p���q�͂���"�� �vW��)˹9`R2m��B`j0���8Y����Z'��:}6�bX�!.?��Fk#邬����!f���SHi�n�HϽ[�4��vA���X�K0Ł��#9�i(��=��:g�?��{�=����Pq,^���%�T��E]�~T��ι3cG��ݲ��-[0�j�z����M���|Ǽ���Ѓ���qpM�]��v��@$s�����Gɒꦇ\C��̂d��>��
9׼<PrQ��o�$�̾�8�$�E|!
jpi>��h��Tes=�s��R�
W�;�?�VM��҄��i��j�;���p��֑�^�qӳ�ʅ|LʑPG6kt���9����r��@C�O�������#�`AUM"#8����҇�!�zo��n{$��=�SeK�4a݇�Ԑ�{Iv�aC� 1,0��D�i�)�ղ���/+�",��-tJ�y���\12�M/���t��oǠ����&B�w���%�"�}
hW��ؚ� H�w&���r���4�,��~�a�N�w0�:��� ��7ǭk������Ԥ�	���F�T��j��
(��i<�8�J.V^a4`��� ��.&!U�}�'�S�~�c�^~1�(#WIFp�>�!�����u��$��/����^��q�^�b7\�QN{����,�}ƈ��q(��2�=9��[�uY�d��|>폚L!wO���$��^�ɷ��gh]^VrX�%EyƧ�,�������2�w��H���<��+��~�
�i�r���9۳3��$�G�I�쬬��I�`���lR���}\�sH��!���m��^���݇$�c94���q���B��@����)�w�E����<�	r4q���VC&��)�iZN���� �|�h��,���G~�\�#ʾ:��ɑk?a9=��v�0��"O�B��)]�g���~�Ƥ�>V�<�C�˱R�`(�=�C}�h���}t�4l8��LT�ɔ�uȞJ�)�� W�L0�/Ne��D�jbw�#�b]ޒ8���}��Um�5�+�z���IH�V#���LH7���\>c>{��GcX��q���8�	W�9�O��^���&|HWF����)1�uN�y]����{�]�8;�p�L�2�ք��^{)�=��.w��r�M����1ZI57;�y-R�Hx���"�X:u�tcf���EȔ��~�mu���� >�[RLh,�5�4�F��f�V��3����K���@Z���)�WG-�	JS�
��w������HȄ�~S���Vɽp(ւ ��*v�
3�-s������`�Y�u���XL���-R�)�U��mA.��_Nއ�kK`<e�je��C� L��K�|0��������{g�%*i�0��h����wcb�0<}�W���z'�$YR�<�Ձs�*�9߬�@��nݜ��d���
��A��&�������'��jQw���|,�t5��5وs���^�����D$�Rkȼt��1#�����o} ��	���q�ΖjKc}���k�̠�UF�u	Shؠ^���4�2�}��֙.�(w���W�p�o ��^h�-�Eo\5'.�v�>��g�ծ��p8��?�)kmr���w��u���3eQB����J�5�b��[�eQ���\`�3,��� Z� �9����]I���	��$<���V���@W��o{�'V�*�}�]����\���q�P��N2��P߁;2�!ujoN���`'bc�~��Z��zi�( O%@-a���T�!t�%}���Vm'�t]��%��RY�'m������C5�[_�=�"����1��D��zO���O�ZXuvנ�сb5��S3�|�����{P�O���' Phh�R��9�����q�.RW�cd#]5^N��u��3tK���r u틦GL���r\��V�>����YO���� �ј�&�&��hXa�9���+�P�1/��&�@�D[>�TMv�RA�ܽe�1�Q����ZoM�_p���k.sK�A�6�gL?Ἕv�ĝ������|�����9�?5�	��D,�g�z�vW@��������a�ew�zR a@���@F�/{ݴǷ�1�m#�S�i�z��.��Z�(k��4���R�w�0!)-|��"@n��W��+��AH*{�ۖ$n.VQ;cM>eԃ��=��o!�I���ǏR�|a�8��&�/ 4`��׿k����6s�p!��k-�HܘZ�7����-�^������3�����Ÿ)�S����I^�1�CR47����F��I�맥0y_WEVe��F��7��1fò4sOEux���h8���"f q��A��g��_��;+XK7�@����6�~}?���o7io�A���W�s�Eq�fM�Z��vO=��$c�FõN�ȡ9�&R��x[��� xl<�]�-,){�[Ȃ���)���A1��"��Je�a�Ƙ�DE�&�-r�Sei���՛�Z��P��vL*牦 �Ц��|�	)_��s#:34I�0B�[�H���6��G�+\|���L[QIbJ�{���J�͓qG$������ۄ�v��.��׳~�GJ���?���w.��:�[�{���	�w����XM\dy�C�O��H-��IRr����C��1�Ɗ�̋a��6{[�(0��ͽ�8��λ�^�-�L|t��-z�;�-B�RgX�`%J��P��1x붯�{e]�=Wf�6�V���O6�S�Č��	Ϋ�`z�#�&F��9��P3�
Y���`��[Tz*���{�ќL�h����Uث�>K~��x�L�P �^sl�%P�C�J��X%�,GB�����s;��]��W�޲�xd�� ���#��T5w�m��6� N�A��݋����)Y6*x_d�h�'���f���1P��I��L��;�hdg��ֵ7뷳@���6�3�����rUU���7�<l}��et���3'�sG��[��"�5�z�����M��:c���cg�� J����HՎ��_�V1䰋�*9��3r���V�ECL\��T�E��,���tr�AG�پ'_���j.�{~y�����&ڥĀ����d�9���FUW��c�	.S�sT�'+�π�Sq��TY��:�n8�_BqZI_XǸ����p�yH犓��*�Q1?|#L�DC�b�6���2�D��5sVa,ꃾ~���xÊ����h�OC�&��x�ͮ��f���ڜ��6��cf��y\�ڢ͐s��zb4#�ƺ��)��������L߸Y�x��"���Q�^>wj�8�x�G�<��^S)������p�\��^�s�C��3Y�	� _+������#K�a�����ep6����<�}��A頊���"걫���^[i������;��O�E�&&r���_�]?ş�3k�F�cUR�f��נFq��,<����Ŭ�BbMQ��!E�m:'�9v�v_"�8��=\W�񜧈��(������1s�@z�2�eN����*���5���^t���b���og3-i����Z��WD�H��ǈ@q1S�'� �0e_��̒���
�ֿs�#�A4{��b�8��A���(,c�?mCQyg�g�!�V����ꎄ���i��ؑ"��:ď�丛�m�zV�z��Ԩ��Ņ�[$����z�%��T�J����D�>�Y��,�0���TWA�y{5V�,-�W�*���Dj5��(�
B�~��Q���2��AO�-�M\�����/�/X1��P�.���V{"�� �;�����Gc�]^�C��b���l��FԚ���Wk&!�b��G�.V�_23�ٕϒr����GS�4����HM{غ��NlI0������`�X H-����.7ra�Y��zs��b�հSy�*�19��3�o�gV�w.9X	�R\�#��A,�F>��4g&�>dj�TA�)m7Hȫ���ŤQ�OՅ�o�E�f*�$��t��iA#�,�v�N����Pj?HYø����E+٧x�?8��_��4��j�t�tf�92rq8��qXV���s(�i�B�	�����Ҽh��^C:5�I��	�mi�PYUJb�f|��)@�)p�|�31ۆ���_���x���Tł����~�eլ�|�u�7Y���ܚ��챧œ��tf���S��*��o��T*��Sto�l�8�oHt�u �|�X�ǈ�R$�1uՁ���_�:�a`��E�K!(�v<|RB;�R��,M���?�!ǂ&�a?�n%������tTf�cݹ5�&����An�m@Z�)8I8���ӳ{0af�'��f>#��F3��;̷9��B�=!����XO��V"�Tރ{��1�z�z̉�!RO�l��n�n�c�^t�p�-:}0�����������۰[*=~�rS5���0M��`�+oJ����-�~�#�S���!wT,��).���J���G��}KX&-�hR���������AT<~)%��~7��bk�D~j� {>a�dD��ld��c�"����t�Y͖9Lo7�kg�ў�M���`�>��r�Ne8o+�xz�7u��Iv@e�V|	�B �D����-�Zi'L�Ϟu���V���,T~+?�S�Ն�zrSz�99_Mu�WN�����jn*�Ґ�S�!!_ �eԸ�d�����>I���rkk ����bI���{�O�gL�����b0?���q�����"�{Z>o�Sh}��x����뎔�Լ�`0����U sჭ
�w�{����+3d/�~�C���pTI�H��HSu0^���	&G�wj��$�2`�V[��?F^J�r����s�,*��g����3V�Sء��ǝ�n��):ĺ7�/,��T�#;�RUq��J��4����+�ڂ�Z�cH�RǷ����((D�]�c�<%V2�i�A��®r2����FN� à�h���O�Z(�}���*��M��g�U������x�4e`#y�����)��`.v�ˋ!)���ܘ������^�(W�hk�>Q�@�g���T�Ì[�B�x�����w5Wp��e�伧�����ƹӽS<6�)3�U�^�@=n���2$�1��G"	�{��m26CK��1�8�y�z�raD�5FX�2�D��W���H�$�{"i��ۮ��,���{�'��o�0���E��l�Sy��{Ymۺi�����x���{T�w����k��>���Ԣ�A(柾e�� �G?��m��-^��gC�%Z����N��LEcL	�8 �l\yj�vE@��7���ZP��BT�sΩ�8�����;trsv��la�P��%�?���ōF��H��X)��J�k�}W'����F� D} ��;��`��T5�T%h�N�0��$��m;4+�p���՜�����{�`��qi�V��BB�b���6ʒ���v��&Y�ܳ�䩓7�ďm�[.
b�+�fP��[�M+^D�KSi�dY�y�_8.x�STӂ�ׁ��x:�ze������)�/�09��?oE��+�~�������O�u94��Qj�7h��V���
�D77�f����ɑ�S��r]Vn�!9j�ig"{��r"�HCd�Mo�
��hF�k�XE8�ԕ� p�~�7�d���bb�ƛ�� N�sȑ�7�C���~I�TO/�d��\�1w�`@�ڍS �:�����'f�������0z�o�^P��4\�Ѡ����R�~4}&"���.�%��:e8�}�ӄ�th�>c��-��?��n�]�n� bGB���X(\��k�X�b���6j5�!؝��ؠ��՟^�T�*�+��/���(��Mw�Q�z���*54޾N���>N�<��S���022�=b����k�1�e`���{̺ۉX�������o6�2yo!$k�a�Ǚ�_�N:뺳�+��-��hdS�6sx[9yL����[�\[����x��;�����͆�����f9=�|��u	.F߆q�g)�$�k9j�������H�2+M���QR�r3���� �8|���Q;�\2r?FmR+�G�.K�l�ܹ5� -�Ԣ��k���B��]�l>�7��<�_^b�N�-6�v��˭�`��p�'���m��S�)nD�� `�<���rQ�G/���}����X�K�	�/3TK�=\��%1F9'́��o�+q����=|��k�y-笕����] Â� �D%��6�a�>W�����o*4`49�܍s2�8B$Q ּ�A�t3��+x��r�+C�γ*����!o��X��\��<ᆀ���`�F�O79�x:~�h���M��"&��ΌkJ�T��X�[�5�k0?F�J<�7�R�<_2�Z2z,SP<���{���Uy��QǰDg/�6}�~�w�gu���	B�R �t���#uBS)��e˳r�dao \� L�%��|���<�?��}��m4�Cz(.+0V��{�^;���~��~�	��6�gE��T���� v���V���D)q�r[��>1��1:#�:wK~ECL��r��Dp_0^��sJu<���S2����XZ|��e�˪��T�UT�Fd��_)��[�'����}	z�{���YA�����ToG�i��^�\Oߡ�R O��hફK"d ���g^5�[�gH�2��l���u7-m�R���@���4�?<���c�$�2G�2a�$ =�3�>���7��7ď�����B^��V9. �}�`���I���*��$����e���e�G��lp	\Ā��!�KKܬQ���ɛ�M��z;��'+�F���>6�D@ъ�y�Z� - �?�`U1-�
�VH/쟺�-��֪i������=�F�����֫Ȟ�RL�gluv�� �J�@C�� J�خ:��@;U֧����"�j���PJ���~)}#�(���"�V���"r_YmI��U�K�]�(�y��?�����B�i���ltN���c�%��� �[8z)߉oj����ja;5<�zoS(�c�m�t蝹Nl�N+)Ĕ��,�!�\�������r�E�=���������� ɉ�^�)E��mږ���U����G�E�к�<W;�^��
��R����f���jZw'ļ����Fr��:�Gn\�|3j���>���2�����W�5�[��u�}�E���>�o�m���ܳǈQ�=�l��'-ZKȻ6ǧf��-����OPlm�Ё�%�HB��2/FX�p�"?��V�tP@������O~t��#8���6ױ30�=h�0ܯ�\>�T�Zْ��?�I�?n6������6�ՅсcP������<;�&��"~2C��3���TMh��̳�_���/�є�����-�[��p/���Y�5ru��"H��N8����f��`��И�d&��>;b��܉��,�.]E
"�WVB,�	�.�gs�O+}VM�l�G�q��^��̅��Co>@�[�AU����m#E�1�b��D��߮m�0ߴ��1��A�MU7 ��LCu�G���x]m��4�����ߨ�:�0�$�B`��$Π�؁p���^d�r�Ʃ��}:��W������9�ĳ�`GR��;,��gȴ9	e��Q�mK�1Y`���p��)�j�a\��60D#Cr���%�w��r��7G��dX�4�[~�4�&�J�_X���� K�*��i�WY�%��O�qX�5mG$l�.MR{��d�����dy�E;y��`=rA�¨g�۩6gCl�6�a���"���C���$�V_�=%�ʚ�Y<G`��w����оS���*A�4�1;�gkF��YW��A�[�Ιm��es���;i32���p����|��^�QYj(/*d 5� �[W��z��N������c�� 2���ݥhA�Ӵ����˟��E�k'H5&����b��Gn?HS'�$Vx����?�]]��ui��v��,��Ll���]I���z^y��N���%Bʰ�MR
V��$f®����(F�O��Qq�@-A��ڻs�a��i������ޫ���[D( s�]'� +��ۓ[F��z��$h-he��rQB�F�xs	%T�\%ӆ���8��Ӆ%(W�萝A�'����VO*&՛S� =��dy�o�|���_"il���Jj�r �:0FG�,�|`ql���M��ObV���̒+;�(�RC^�<�BGܦq��A�GiJ����8K���[��g{.	�kg�UƤ�^B�%�&<AiU��5���r/��v���Gc*A�E��mY�K���+��+T���	
�Z�&����{<)���YHKf@����g��{�Yx ���ˍI_�ş�o��<�[4�R��RM-�z����ʩ�]Ė(}�gI~JnwdX�ep���x�0��6�')�w%xG�wo?+�YH���)��%����d�u��?U��{���vg3���
����F%սю�<T���e��,\�a��a��v,e�t;�w�u�IM�I2�����>��O�;�?[���?�������
�yʗL2`��M��.��J�t�*���p߫��>=&|����F�*�H�2��9um�w�RPtQ��@����Wz�Ѡ�>C��;���j�1͙b��lOB�r�Y�u\|��}r�XrSɻ�:�ٍ9b���J�/�b&ɡ���y��y�Q/�|ְ�.-�����3� ��x���B�n&�՝v����|��I(ߔ��lA�P���\�q�C��dN%8É�I�?s�q]hb�w�=��)�c�ŋ�Ye��� �:��x�_X����R��g��aNK�����D(�w�FI
���~��m=�w (����`��2S  C��ǁb�@ZFԀ�������P��ӎC{5�`5��������^U��cO���hd�*�C���&z	���� ΂�mO[*&�`?��5s� I��d��1�����
�zj`LL�]�� ix�'È�Z�I&�c�;���M�?�"�X�����'�z���:�P��C�� �L��������WѽP-D��]ʾW53�n������ɔ�Ow���j�%�P��eau�E7'�ĕ�5 Ӳ�n�P��6?fˬ7�X0�F���߆(FX�Ϗ�z"����aƾ�!��ʓ�\��+�;E�d[�F*�o�m�Y��qǖ��|��0�����g���(��:�y7���f��4���ǖa�V/�Z`A��?�=��Q�lˎ��!���b�����h�x��z]v%#���N�K���=+�[��(���i��-Ǯ_*��r?v\.MEB�@�Q�ʶ~]�tirX{� )���0��$�>Z&�5L�tѻ"昗Ѿ~���ŃA-ճ��G�N�h��i����&x--D����
��+@�������o1ѦY���ʹ%��|����M��]
T7�M�/잞5�r��Qr�Ҟu%�ٽ{���T��,|�E�w�gϘ��؆�E���w[�-�(*���̈�Sk�ɓ�
:読u� � ���Ƈ����&��z�~�饎e�Gf͜��h,x��)�[��y����!��V,�}�*�ɢ9c�r��jܔ<�`�f��B�*�»�Jʩ-/����hZ���ãH��@rj��%�``�	�
��WI:�$t�B9�m�U�M,��3�}�	J�)�w95A\���@3-�`����Wǜ)��2�����Fִ#�5?<M��8Z� ���U��=��l�����$�Y��_�Dt���Hr�Żr,ğ7�����r��4�NVˌ��3ns��P)֡� �#�R��/͛Jr�\���'b�>�1���jam]�a�����u[���۴�j�y ��7à����6�%��� q��������7�Y9W|d6�v@�ĻYYnx��M:^�n]73(�-�uqR4�b�:*���MƔmUK ��i6J:�,��է�Ί�ǱP`�$)��͠�1�뿪γEm4~T�n�6$Vo}���%� ���F��fȱ]����K�8B���wd��w'����~�_�Cx�_&G"��^��r�������(�ҭ�^���У$���-�o�Z<��E�"��U8�k�w�ؓ�T�$8@L2���[�ە�*�P��"K���eD�2���N���t�X��� (�x��5(�0���3$�*�/�}4M�{��z�i��(�ۈ]g�4���c���f���=`�L~�ā͕�^��V��)V�x�b>���hH>h:�%�P�����'�����{�g��@j���0G��5�<������%y8n���R����?����� k8���M}�j��M}�|�o|���R���Pn:�ʾ zT���[7�� �Gª�x{LɽS#9=�OIx]�B~t�.�$�bz�`����+ҭ� Y�G�y$gaU軝Y�5��T�CJ��쏓>Pe����
P��&U���������)zKKe]���sġ\��I
����k�>xY|�k��R�)�$�oH1�fCT��� y�T� �.�uL[�k�7��;>�L�/�R�^����R�>�Y����\�T5�E�w3�xt�6�Y�c�Ċ�^�Nυ�ma����m�C �O�ѱ��+(�of,U4ކE8�8c�t��J��*&J?^�P��2:���iHb�����졲ޞ��X�)�#^��ȹ������,�� ��g׫���	-JzΧ+ �ŷ�� )4�;�4�n�tl����M^�[u��Ȓ�N�	�����&֠������	Ѯʕڟ�)N�F�����+�O�+����4����lc��\�<��*�i��,��[qP��c"##?<n`-i��[T�
k`FSO} �Ԥ���h0�^�؍]X
�>�E�d(ɞzfL��Ϳ ��Z}yi������l<���S�q����㣀�K��ح�*9����b��a�{o��Zb�Gb�����a>q�&�i'�A�+VnNs���a2~�V���lNq�:�s����Ȩ0��-�P{�@����m
�x7�z ��CK鱿�G'�����i֧}�YK��b�;m���c�e��(˟��J��`<�~R����"�c V\�2t��뱩,����l�UL�vzG��
�k�3��Ĳ<��ciG'�D4���� k�����!rOqy7�PQI�䐌TV��t�DCʹ�s��=�����xq�D���I$�]�^�NFg<���Ӹ\�ci0Ƚ��~���y�AN�D��5
�e�XKfM�7�HE�R)�4	<��{�h���2ʳ�8#�9�<�UcͿ��ba�$c;\� �F�-��ϟ͓�JY���9xS��OVt� -d̢��ƺ��^k��(�XٛH1"�c@@�-��@�Sy+ׄC#�Uk����=*0�@^:���1~�'RZ�՟������B!�E�E�>E{C�m%��t�z��Xk?��6y6Pc=ڣ�$���������1=�T�T��^�����{������X�� !�L����f/��$�?���k�[ߔ�]�b�s0%V���}"�	E-��䡥�c�Z�-�vV*�6�HK��u���~���BbHc�$���W�1���pHua�	o����2)5��yį"l�4�z�gІ�+r�����"o敒+Q��{I8������?h>�%���g�A}o-��q��ك��{�u�����{@&����sv�����%1�B�b��u�fYd�x&5�����&ڐ��w��R��!=�9��)���F�%}��o%�ܟ��LtI�V��G h�yy����݇=%��UI��I8.�ބ5���e�߯o}!J7O�ځ��#���q�?c�4c�K�H�qG��3�����_W�r�؉D[�X!�V�䣋�<>������;_)��mr�rN�_�4���H��T%	8x��/֜�6�`�ȫ޳�!~��5^���9�K �o�k-z������,��L���i��y����7yK���x����!�ZD�]#��v3�CE���)S�N�{����\�
+�U�ZM˰ldo ����oty>�_Zt��Y�{��
)��Z�/�i6�:X�NF6r�U�^��0�k$�I�-���NP_!ը��,��%���
v����D�T��As����?Y��������ˈ�@i}�>F�QᎡ�>(�3n8�z�v��;�#I
�d"� v/�O\�|��F߅XV���%�3�������J*�2�SQ����DJ���
��J�e%��R5�qˉ�<=Bͅ��a/k�xϻ_u �[Kt��H?�	
F�aEz���K�=�eGR%>���r.x}Ҽn�����;��b�-@��o_�p�����W���#�k��#�ތ`�h�85�(����jC'1� �`�;��|q��!���l�Xt�!����H�Ck�b����.\m+ݮ����K��+gi�G�*�9�8��M<W�i��c+�SS��:�5ʍ���<ni��ѣHo��hr6�1⿋�i[���[��q������tȐF�("YE4 �����cU�"t ��a��=�ȌF��w���SX�,Af��zR�1ѭ����oп������8���نER
�W�����٠Y�;7��;k���L��֢��V��I�o�:��y~؍^ߦ��깿�A�T�"��V�צ�3�(Q��&��������R�t0GAa��㇁�&.U�a��lJEp���|$Ë=Z1���~`d|~)]ZZ\��я"�Q� >	�V�z�fKKA��<�g!*6�y]�G�ʡ�(�#P���7�d��z����w���*T!�T8��"N	u���a=�&MX�ߗ��!?f�i��v��~rQ.�Á�t��^̶,(�M�R�f��� ��0ժ^�mJ���Yu�K��uN�m4��S���I;f������O�M�D��nV�m�2���o�:�j#������}�;Bjg'����L������t{i2�XN�nQ�*`�Oq�6��c.G������mi9_���=>�~����m�-(�����}R�;t�|�E��.ȟ�/>#Ћ����l�C�dO 8�����+��F�y[�T�����[�S�<m������׷��s�����D�>pH��$=��z�+鍵�SQ�\��^H]xTugpE�l�[V�S�6�7��lk� ,�?V�8�I����L�>�t��l>��eP��>"8�-Qx�I&�Vn��|ɏ3���ٗ�<���F�ѵ9c��œ�#� �ج�pN����N|��c�6aȋ�`�S�1-j�$�"iO�(#&��G������efp}�h��BD���#���[#�S($��`K��k�j�߮�i{rR䨬��S�6{^�[�{֮�Kt�UX�N�D=q7��b� ,���&ApObbs殏ZB���:���(T*�7,�@�3�O���z�/0I(J�E��s�O�)�A5{4[����	�d�;��7�z}��ʪ6#��S޲.Q���yC-�;$ �ot姠1�u鸢�5d��޾:��}����ƂnvvR��I� gI$>�ώF�-������6�У�R�q�_�`�����7�e���o�վ1D<kx4���E#Z���&��t��q9˱%�
q�ZFX.&>"\��=&5�֒�-�a�g�SR��o�h�����9����o�q��v�l{��E���HԡT�ac�/�Bܪ�6�ۮU\�j�;|{ߝ�YwyԥW�e.N���'�]=V�����B{.J阆��zG�w��8�h}D3K��ac>pf����E7���X��.O���6�����VP�z�����1S�YAmSË����O5�U8n��h��C���'�;2OŨV�js�q�@A)�fJi�c�Y��Y�j�̡ܢ�f	��aa�,�&�\vk��³!Ws*�fK����_N���!Î��"LDN3m/��O6AQ���,���%4@Z�"��FO��o櫮YC/�j��ZO��{�P�]��#�ۃ�v����%���/��_W��J�9�$ͷ�y*�V�#�	��mDE�^:��Б���ǔP�zR���֭n���\�ż����!c��rv�����
 ��^+�yd9���/{&��=<��5v5��e���>7�o�����:˂��h����s7���Eg���6��%�>)^�Z�Ǧ�ę�c�;.a���Ej��?�٬s��Ҋ�>a�;vXJ]t2a��c�+�X�EH��T�e��.�ϊf72u˵�	Ъ��&`=#�Rw����,K��o9��֟��PR�8��ª�B�P!t���߶O��7m6� �ف�鎵Q^��^Z6y�|��Q����r��&�����6����&r\�b@�Р$�I�A/��c��� DI)�D9����zj m-�e*-b��F�" �8L�E�\ ���5W����f�c�Xd���ng�
s�Q���� |��
ӻ�*,a�J	ڈ��$X(�K&����n�tf�����Z�����Q�zdZe��a���4�GU2R1���Ik�c���@�����q��1,=�
IbH��W��Y[�y:��F$mg[��%V�]L�ɶ<�\O0?G:���3q�\t�Ɛs$�d�F�-s�$�ZĬ��4���B���<��d�k�&G��Eܑ�9�������������j7��ݢ��tJHj�l�M6u�Wl��~^X����U�-]#xO�����t�{a$�ͣ�D��<�0���d��@��w�BI�^r�F�c���F���$�m��$IM�st����jN r�������%�s#�񳛙y7�C��C�}��ܸ�����.l~`Ԡ(��7���6��][`oh;�~̞i��G>�#U�	V.��##���U�g��=6^�6?����7b8��"�a��C .@
m�לx���:
ip/�T����\�\��@6���,�u�c�4��ܩ��"��Ww��ˬ����XR��׷ƵpN(���ӄ��F�����՞>��m��ȭ_�װV�-���r�z@�g�x�R�5O�ʱÏ��5h���/��K�j���R�~ʈ�p�
������\�d��1U���>:S("�{$䑭R>(Ip.�kt8��8iz+�fq|���`M<Ju�P���y��y�#���JNI�G�7��t���G��i��U'��9�$���А�)�iO�0�cm4iM�y��U:p�k�����Q������>��߀��T��t٩�c��Q�VyVkmF���n�$�`8��N8���h��N�h{����rC�����0GǺǼ���R _��~M��D�?��l��.�3���q�	�k��}������C�ƒRpB���PD �<�ю�u�RG�����[d^�b<,���>�i�(���A^�`b!5}�q��O����/)�5~��h�G���!��,�PPXt}`}�4p��S`WQA���b�� !sّ�M��،�Z�dx����]����ZT�(i�g9��y��<�J��yɪOQs���m�=��?@��n<�W�_O���[�Y�&Vx��I�Gt#���1T":�/�T1��j?�qH|`���ؕ;��_b�Yl"o8w�{�~&��Ы"rGէC��
���V����/;fj�M��>��U-F��h�MI��7���v�q�L�o��٭�E��?���<�5�D(19��Q6 e�[���D^�A�NK�^ݚ֫����-T;�/�;�PM�]�ʶVO���� ���Ro��Uhi>c�q|4B��&Mұ��&���8ɀ]�S�ˑ$�ΰM�H
|Ʉ3/☋���ޖZ�ۤ?�0�����k0k�Fԉ �l�̆s")��4�Ǟ9bNy�\`����a���U1.��ACNPެ!+���Kh�y����/�%0^�,[3m��%LX# Hy��Z|>M�%�Ē3��a�!<�-A-UFCz�ڧ>&���20�`) H�x6Gcu�22{d��wq�6y��mbd%�N��t��8{�&$��b�*o*u�kj�����t��[x]�d�]B�Q���띚Є��	�;����G���`�������ȄĶ�[�xN`Ξ��_���/�+ :�����̣��PLE�J(/� �	 ������p�w#>7��g��4�� �KU�
sx��8���-&�X�yҸ|�7�.��r�Z���Ob�9���%oq�rO\\b�Oe����O��Ag6I����\/\s+�g�f1?^VX��wː,	���D�2d�_��Y^��[T*?�/�_<��ŀ�|W����Q���1�a�����K�>�*w��FU�g���1�K��M���	^����Dy='}9��h&&���tOٙl�=?_�ƪ���p�ϕ�i��k�h1�W�P�Z�m4��&K,:�s���ؐ�00�ق�7NW7�qK�#ˠY�����T��IV.�|df[�ܲ�j�ъ-�:�<��WX��`8{�C���zs4����P�v�X���;�q �Rs#(�6p�1�m��HO��F�w�9�Č�ϪD�\�'3�C�䬠��\�Y�г�F"�FcB�]�CGTS�cgŏ��`?�-A]J%�'N�uw�7�ai��	4`�"��Q)AƱ��,_�	��$��!�c���FYH�R`�lh]��˥���BK�a"I�jڎ>q�NU��ԯ��-<������AQ�����8� ��p��W�԰��A�c\��:���(��,~K0�0ee������Ǳ��f.W��$>c������`Q��β`y1�zO��.hƂ��e�1�3^&yv��4]�/&�*4�<o�^�ٺ�S,e�/�%�m>Q�wDax�򪱭%U*��^�� ���p�E��v�\ �΂w,��ӛz'���1�u�|h`��s�O�Ad&Y��>w�"��
 s��@�ʤ\�L��#Td�x�#�����GJ��n<�!5l��|�B
�L;ٝM"Oņ�6�E����*�jh/v�S�	C�8�j�hnS��zĽe;�;���|��`�j����W3x�*b����L��Yu�Hy6I�i-iEJ����ktma?�k<�M��yD��T�îDm�&@��"s��٧��M}"�5i�QH�����/˜H �;�`U�C�}J��f,e��*R<�a�ܦ��Y�^��?-�Gt�BW
�) CZS��h>�[R?lzRȱ��(M� �t�"o��͡d]���&�-)g,��׌���Envi�SU,fd�+Y��m͜Q��\/�6G�=�eS�QGB;{��qָ���F(8�wJ#p	A�\�z�Q-s�\( }�����Cz�AuvXWS�>u����~n��
{���Vo���i��4�uVP�Z����lk;����:_%�Ӣu_m�O�y��w�j�*���[P>�'s�y�$��P900{�uw�*�d��8A�@�H����ǃ�>|�Z7i��ĝ���M@iD_� �A��4��v.���sA)�Xl�O��	`7�~�/0�߫�:���PA���25����s�k�m�&���i��ˢ�F�>z?��v��@�⚉��,��@�Qd���X�n�t���Rk�k"� @!F? m�z�z�{m��P����u8�p�ōk	l_p5}����6�7�w�#����F����-.�3��[�CR�G=��3w��@�ߚm�MgUJ�<�Ks���b��$�6�����-v�֟��7|}?C�Nt`�6?娭�mrZ�mo��d�At����V�Uaۆ�b������w�Ԙ"�ŷ��bW:)����uZl�i�@eߵ����u��O
�`�k<륹���������,Z8ty���A-}�� ���'�a�t�����n�IMjNlɔ���@����F 7��03�[p�5���f��w�����i�&�J�y��{��S��P�U�|.uqi^H�Ƙ|���]�Z���-)������x����(MP�w�lմ�AR@��5�by��mku��g-Ī�6�䩁۫8Gw�P����@���Pl7�.��8�8���5AhXvdzt�Q���vQ�l؟���pTz��0�.�}$�O�r�����,��D�r����`+d���'1+�8-�N�}Z蚴kg#�y~A
L4	�R���X�0���-���>����3M'A�ʸև]k�NB�P�Yg���]�^C�NB1��G5�j�^�~�2�Q^�$j����NW)G�~�z�셿[̮��ix�R���wxC�b��)��@�FE��Ã����mu̔ڪ]�bˌ<�1ԑ(���̮���c�1�VE����^�bj�	+l���.�/�7�R�l8�~v*�[�T�y3��.X"f]�#1���5�@��H3��Y�}(��2v ��`=��{qh�����=�ڑO�#F]����kj�E
l}��W��Lh��%�G��2G톑Ų��(=d����k\��.�\A-�'�>![bo+�	?m�QꙉA�����l��9�1ϓEH��D/6uۼ�1)y���8�xU�}�ug3����DO'���̈�d��H)��|�#	/�_���tQ�)U3��1`E�f���G����ܩR�~�����"U�3 xI�"�/����ݒ�@aR��h�H��6pCdC�w���Zt��SU��dx*��D:�3�P^��/�v�Bm�� hJS��(o�,��G�h�����_A��L��>�;^��˾�2�����l��(m���:%����Ǐ?����~�w�,'��|�~�t��z��
�ɎމZ<h�:�e"��+��k~౨y����}/����+�r^��C/@�U-�	�����x-�q���:c��N������;??���-�H>��q���
�c��:afHd�zl`}g������T����|,�bx1:��軸��`C���lOh�C �� �4����LL��!`5r]��,�J��ݢ���W�pXѬ���3Tj���	ʇ�qH���L��qx�W>��5�==�e�?��,^���8&���u���C jx����M������E�
��"��PKH)}�>2m��O:�1�TX�/��I'���a���yf�C������IC���)��ʴm�U(�>̀*\Zg�#���ER���(� �4<lZ�/�Hu�2�a��^	=9����C�e"��o~��]�B�jh ���	uR�\����]�3{�ⷊ��b��+�J`%�Fw��Pf���#��l���v�87i�.B�S|*���#��A�`&5�>a�Onc���x�R�uSx�7��>7q�;;Vk��A����k'ʟ����]�+ )�(R'>;V���A.�S$��^�I�9�sۛ�l�vh��Fr�$�ta��@�i`ӧ/:�jQ���]��C%�]�h�h�=���qV��'G��a���V�6D�Q�t��d��G���'�
H���6��ǁ�Q�U0舞IJ0ңgC�y��2 m�gT��e�FupAE�oG��M����!@�u���i��6���ˈ?�NޘC���z)�l�P�0<�����Ɓ�]r*��$�(�l�w~պ�|JJ��{�䂕9Յ֍��#S����ύ`{ M���y���)�|�À	� Mث������>sB���R�_��tBf)-}�ٳ��;+��,���--T�#�R�n/����
yU��˺��#T�^q��D�X��8��� ����S��(V3r�������@V�gY
T�#����H'	��|P[Zc�ʺ�ߜ�b�^J���E)�s���bt�"��U�[�e0�h9�&\���n������k�Պy��d9���V���A��E��h������p��N��ž6_M����1,��+��.Yb� �P'���K���\�칁q�esoޭ
�X5�Q�Q���9��ߐ��ǜ_cEl(7�6�Zŭp��ue��m0��(���Dk�q<[��V*8�����tu�8�ĉ��\�@�/�.F���Ku�i��["��~�� `Pn?�p���w���y�О���*�����o�<.:m�v
����t/��+_=@}ե�/M:C��y����y��F/T��v.���T�Q1�AL#̍j��������c�;�ە��%>@	���Sܾ��C|v�X�B��&�lk��(S��Ey]��A�/�-����pL�R���u�;�#�.��� :f�)�/"
 ���Q�1-?w�>�?U2����İ�!��(�5<Ǟ�֗�S�攒֭�:�Ӓ�:�3�枸�ȲiIt�z�R_��v�u��>.�#�7g��$EI�k@�T�YT�M�f0�&��^D�'�w��?,D��09:��n�{�B���_y�n?j4��*�H�ͩ����΋�g�F@-�a.�s�F��[]w�Ǔ6U���F|@!-��y4FY�&#��=�񁢦�j��d�++&���e7*�1������߿���'ܣ�&�*�N ZCqd	[G��5s��M���rM�~`K`/v��j��(!�����a������4��*��w�� �/$������0Kb��!�åj��!k�q�>���BA��x��&��`�^�VgR�0*d�Ɯ+١q�Zy��+b�ixbd�ͮ��͘��E ���l�<�_��ߍa�W��ꨫDU+d����c7̤���{�~_�\&�s.]�֧j�m���.G��Ey�?��n���y��)?f`)p��}���c��;�� :�R,��i���g{��b<��3q%L<���D�~d�r0���I~�4t���Q�q���z$̠M��Z���]��t���<�y�7��7]�.@o�f��<6.ԋ+���s�P�)�V���E51X�pk^�W� �j�LJc��o#��_�D����
s�׾{%�,[�N����i�5k�y�)|���]��_d�[' �� �������t��蝀�B��E�aMxAx(�?i]B8��¸>���!��X�j(���;c�8N_Y��㶒"�Y�>��=l2+�89�?�)��p|֒�S�Q�Zw@jL_�ٚ.2?�.�aN��9<�]�e�`�|�&�G����ykt��n�Y���E��ϑ�oE'���u��k�Ɲ4��c9�%%<���v���W^r��0k�~?���6~m��]$���j��&��(�f�R��#��~�����C��J�&Wk9�4qωt�RSn�[_�MF��T���.#y�B��r�5��P��c��HRӎ3{�!������w,ϐ�٘�#.�� Rj�w�\ ��F�`h��p�`�hËzPS��y���=��f��)T$1ܓڊ�E8���;.���e:�ozΑצ���B�+�"'��.(�?u�\���lj�Z��ˁ�F���#G��;�^�8���J��R�<��ǟ0R��UH59�����~8����6���s��$���՚��k\��?���z���c*	����6�l���֝���כ�I|hf��A�y\j���G���7�i��$@��K�qm��-�e�:t�o)��?�q���>#?���a_�b�B��A���@T·�&@+W�ɒԖ�(քxN^L�m�ߩ�b��-(����2�����0�^Zn뢰2�̮;(�uD4HjZLQ?�5�x���њ�.��~�n��[�2]�Y'�4_t�o�UC�Oa)|#�+6�^���Jϓ���G�F�m�t� �΅�m�t�+��m�G�\3\�&�S�:�)��k����`{`�y�g|Z�U/��;Cw. ��Ei��̜�@�K7 �-�� ����`	!�	f�f���&Hv��l �x�p���E.���>\eu�U>f{w�IM����$N�W�S�V�e��
|����-t��Ⱉ��bѪ�����L*(�)G� +�<p�Z,0���i�E1��3u���\���O�(�*��zV�������?cst��|9&3l���[�n׫�{&��eNz�*�F�l�\sp���������;�78��Q2��h��ou�(!����lZ�������Qi��a����]!�Dɉ�p[�k����h�Q�i�s�|�ya~��i�Uy�����ºr��^�Y��ϊ�N���GiL	�4W�S]�Tg�$�@�:��i�=�j6����X4h��c\�˱�̉M���#A��a'8��z����#[�i|N���U%�AD�=O��76��A��WW�ؿ��]E�z��(��o�{Ios���6KHnBf�"�I��܎�7�	O^��Ys#�����<�C�t״���f��!+�������ճ�X��1�x9�ˮ��aZ�.��?_�2�^�M�'Ӷ-H����hA��;N&Hs�s�~���B�E#[�߹��d-C�	 Sl�+�6�p�U,�#߻��4�7z�G�vw刚[�X$#�j���5+%�ZKI2���Ί���/i��'(%Q��=��E:���2g���xp��²�Zd�K��*���q���k,Nt-��=�a�g�}�c�>�nՂKx���e�#8�lr��RנoL��\�^� ��|�WCެ0
��S�hX��r�@��W�?_
�*�,8�E�a吳q��M���Ǥ�Uh����K�hx�ڷ��!�����$X����0�q�c?Hȷ��	���,6���ɵe��9��-��d�t�1㏭��E�'8:��z,v��c1R��i��D]��ˎH�� ���������i\
�U�,��p5��ie��HZX�<�q^s73Q��l~F�w�6��U��Xs�1w����~�c�����\%K�����h�����.���Nw=�0Ɲ~4-t�/�?T��^�/B���@�LP)��&�$��f	����jo��"C0�\��~�s�z��6"rf)��B�O�"�D�5�9I3��ѷ��K�<����>g�="]?u���D�#��#"~������/�~��os<��,�d,6rT�k�{�� ���S�>*^C�H.���F3 ��ƀ�]�W��a�7�5�Q�uG�(K�^�6<� d|A�[lvS{ʆ�E`�b��7��θc�&�#y Dg�>�9�+|�]mqu��}�� � �]�F6����rQ�b��oj
�""Fq ܈i�T��xJ2B��<:V�*����(A?��
�b����<xpDlR�j֪W��������g=k��Q4.e-w�<������'�qr�4�t��3C�%}=b5P��o�\��W�C��=�|�6�c\��n����BNcU��	�g((*Ί����\�o,��HN�̓������j�������]�D��ŬڐPN{?�'�^��F�$0��<���ȣ��C�a��8d9:3,:�~�7c�U�Ak�2 �9+��Q������~}��*��6�Z.t�N+r�&=Vxw|{�[���TZ�t�D�?ƂR�DJu����U�!��۰�F�]tq;��s�3�5�|3�����|ce��Z�z�S��m����J?���b��޷T�|.��j�3NȜ�Du���׽c�.�8|�ڥ.Ӳ�}xG*���R6��n+����7�5� �8}<��z�ʘr��?$7�Ԩ?]P]�����̟^������$Bx�E{8á��0���p-JR�x��%����*�c�!!$�<��Ds%3a��I6�0Ff�,���eJJN��&�����/����	�ía����|Z���H~x��ޓ��WB�����*�����݁�8� e�G�K!
YZg�I��1����ہ�e#������Y#�'������ ���e�դ� :�k^�4��{�L������F�N�p�nS��R����TG��:��ƃBG�0�S���Dh�ٟ�I^���K�tߠ����VԋP�Ŝs2%9�ܻ0�|��ٮ�ISX�����Ֆ�
أ��3��/�-��g�6�!hT��!J{,Dw2�{hc�Q'�^�߁>���ם$M�6_��X<!
6W
yu�X� j�	�X�>�v�3oo�b�^=�����ˬ}FND�P>�I�q����a��7�
�ȃ����W�N.�|�])_5��uQš�o���Yզ���$gw�YQT��B��Y\F��^�1Qc	���6{�E�T�=o4fF����@9z���:��S�p�;�q�̌-!2%ĬJ�-B�x~�I�D�
x����y�bQ!a��4�}S����)�R<#E��U3�$��r���/TT�� �	qhN)RFi�ml$�I��l`�k�R:��e���>z�@*]၃�E��_�[v����&�R�z(W�cS��&,��?��v����.;>�ܴ(,�3\��29v~1����|��yiU:�[|�l�	��e��L�6�I��F�yw��Ք�M;I���j�^�D	-����V�nL�i�@��"c�,��:T��Υ�:�u�>��̮�� U��qW��t<���9����)�}�U���b5]����{Mh�~g�2r�H� >��i�o?�B����3v�W���~t-�I���q�����P?�6K;��o�.���I��(�*��M��=��j�m��a�87o_qh�ޭPk��{[7I�ѵjM4� $Q$!SL�^;�Q��w `��]3.��Z6��|P�"�^ ��^"���6���'Q�3��Xb|is�G�6�����u�Y���W[�m|�i^��89�]s����4�e�4��PwX�d�㿥�g�A�f����7�jvۚ�)��}"������[��3��i�M^�YCs����F��ܥzi�E\�YJ+����g��C)�3h˜��e�F�l��/�5[!�4�΋<�෾�J!�� Ң��547Z���SZ����`��������k��/�����|Ix��fډ8S��=a>�z\�DEcN�s�E���q���d~?�Go�A�e��$S��d������3f���4:Rr�͡m�P��9w�@�)Wx��#��^�0�]��<W�0��GI�jt���Z�2�cJǫ�)�l b����DV�a�Q�wM���fW�� 7bߵXo.�鲞�l����j9�yg�Zʚu��J���y�X4�!uK��p�.��$~�p9 �kT��f������/�}:��K��߄>+�`���톭�@�%���b���\��߶��n�$��7�I��`�i8`�׈���B�����@���Gk ׃d�a+�e"0�H�B�↗�|BY��0�'8�J���[na���a@�nK�?"�M�qf���ܣ�`���8��J�I���-�����n�%����Z��Gs�`3�C�0��7���݄�<�x0�g��kzU�a����0se5��H�YIk���=.�r��J&5�*�K0_έ���VX��J��(��g�C k��c��v��=�{�|������ZŮݘ��f���%*�Z�A�6*���]��j/��4/�*WwIdAF�Ϊ��[����y�M��KQ:hl�����ӧ`+W e��|�.�$��c��y��ռ' CBa�h���B��Z������QB��pψA�|*�x&i��~�����x���%Uq� ~6A_)Xv���D�x1�҅D+E�B�c|��8	���=�e?�|��O��b�OyGK='*����ԥ��S�\>a���e���ic�֚�\[=~�#�H�
S�ѸJ߄Я����I
��	� (]G����L�D���/���3�ӗA�9��z��m��!�L��m��Oh�|'T}h��c�_l��U��рz�&��z�\W��B;Hk_<�􀥤�\�����3��,P��@>��)�n�Sk��6�ɺ�xa��Ih���>
�B�9*����:Դ���Eae��^ۼtC���0���X*�����A9A���^�}��f�}V댌��=�s|\"�h��+`+�iPQ6�]� �
����� :��Ę�jn���4��[[����6\M�=]Wԥf2/�)��<�RT��TEXG�!VA�R�*:P�_磂TǶ���JLz�o}a�d�@�,%��P��w��/����(��4����?@��|%���*�z�ʐ���G��efUU[��� �b̓�,D�BZ�C�ي;�nǌQ��E~��,������jH0q~=������<�%��I�Ys��Ƞ�n��19O1��߽L���ҕ_�۪4�V�(\q`'����?sŖؤ�P`Q���%���_4���Z��nF�'�s����Y�R4ǀ}w��L#����ɣbVI鈤t�EA&�;(ގ�J��LqB�u~���)����@u�9���0��Jd�`�9$����iu�V����t���_�pc���9tT�/��K�GW���4�n��l;��Kj"��7��?�'=<dx�m=�g���[l��奉�|��HL�b*��TE�D�ֈB���M�������X���Gx�Q�@d�X�wY��π��$��tIՔ�!�	�f�ql�)���re�n�b뭼�U,�S�iz��A��m��'� �9�}U+�/�p[�4Dy����[{��&�d�,C���?�4U�Ibb4 ���:�o�Yۦ)��x�a�a0�W��<@��Ե��woN��n�J@�	���4�;�6.	v�i�����H����+poNd,�ih��d#�%�f�}2^ Zx�"�Ӷ���{�m�7����o|��/�S輭��Q�C�i?Ƣ�.�z���{�l��1a%���0�!����r�S�8~�x���_|�3&v������X�c7M.�#���zn�G����nr.��c�@���������~*��Y���-����|�G����k�8tuG��.lBxqi7��W`'�k�ʚ^�߭�F�<vV"A%�7;�=��%��̒wG x�Ņ@��h�sjZӖ8	�K8����_1�$��������_�7��v�mΒs��[�+I=���l�޼����-�;V�� ��8��4x�V7|��Z/�8�$��/����]7���Y��q�q(b���p���*��h����&�4p�V�S"��#�enM���r�,�w355�n,���G����wX>0VD�i��ʎ�����Mܭ`3���´��f̿�s"�@�u��$�����EW�<\���o��/P���VŲ J�ē��iM=r�ݔ���5a5�Ѻ��x�۰���wb?��<H���P��Ӻ�V�u��@qۋ��;���q��UȪ
��v�\��ŉ�Z�|�|:�>Թ�UՊ۵1����O�����(5�mPbH5�q[�K�dQ�̀� �T���sk?����o�ރ�U����L u��+TC�����h���-�o�fFm(t6�kV斮a���+\�����^�v��	5��w�s'����M�e��B�d���Rȷ��/TCz �^���DC0���<�2�k;b=��1-.���14k#Т�j��Ƞ�ߺ`�H�ʞ,pz�t���א��U+ոuC&-���,���fӆ�˭��:�Ӆ/���lcTb�l��0{��vi��K�����5힧o	̬XiZ�h����i���mY���o�4�}֔��z�)rF�:Q��mC�����u��ɽ+
}�lζE�˛u�/�"M�9�t)BN�Ǧ]�$�s��n�m���ŋ��� �݇�ʁ�j��7"��N��\Y�b�G�(�����;~�;����,��� /�9�:F��nn�w0�N;#�u�d������ͦ�)U�#�m���t�)��h:�KLo�PP_Eoc��t��!>+ �:^md�*�Wm�� w�@�Sa���9S��Xڎ�Z������ZUh�\�"� J��bEn� ���>��&Bl�a�3��JD?[?�����+�[t�]�H73N�bI�(c�|iط�2x�U��G�zi,~�dMTi��\oX�诘���CÐ����S�怴�|ܷ�h���%�Үw`�,��h(&�	s3�����d�	�Q�nS�Fn��v��P�����d__�S�bO�����m��u��Y�sO�ҕ/�j,�in?.�_ѝS��h������l�ZE�Z��T.�s�t0���*�s;SD�ByD)�+y+�%Q,�k�H:A��U0�Ǯ�5D_+��sn�����tpC��TT�v��h���~f���#����n�[ݿ.Wl_�����Uu��L�X�Eڷ��R���Sl���|Ѽ�۬���I��T�2І{��e�4K�g+�RT$��s{����Ј�(<�6�ӳ��M��nk����M��b�_H��sD�PRR�gT~0ľ�!����c�����t7N����ۧ���
G����{��g��J[X�I�����A�[�
::rV�^����(���4U���5�K��e�B�@<�����h͝'^��!�
�~`g�4���g������U��g�Y�r8SIY�3i��p,������j������wkɨ]|N~�m����i�J�0"0P�y�h�`�f���v�j�3�P����Q��pe�$)��/�R�ܸq�"X��	�=�S�gHQ9�5ܣ����=��G]�u�\Լ�~���;��6��1�m�X|�=�ߖ^C�_����1�o��3M*�����Q�+v����|�bO�#�x�7tF��*�v>dZŋu\�����/�Kc�.9���W����TQa�o�&�*�	�l���P���ZV�J(����]6�Hb�f�aS9�`�.V�ɋ�G[<�D���XHd�k7w��9���(,��\�ug�@=)r����T��<�Å��f�&&�^M;볆�����t;�!-����D�������'�����]�lA�`����/V,�׸��
E16������� ��4����	d(���E/�L&{�a���RL����U4m}��?%������B�r��=|�����,����Z=��5e��6����(2��hy�c\�UQ�؁e��ㆾ.!^{��G�?\h�\�Z���Z|�<�W�X�4��9�T��1�\o���T�@���� ���h�9����Rk��1
�lk+>�o�@o�Z��Ȋ�Q�(�d�z��Zv�(�B��l"|�7>��yp��� JY�,Y�@<��y~j�Eޓh�cؠ�D'%1�8)W9��#�9m��/>�أ�ŵJ��Zv��Hv���$���D�$�Ќ@��F��,w�sP^���)k۟�_�z��0v���n~���)d�	��z�#4pQ�<j��1���gFQ^�j�C=��d��<�φK
kH��[�u=�rJ�*&���ez=�݉H�Ȅy"��X4}��Ma?��%�R@�����0�B��y������g6b�1�ժ �FG��@����ĸշ��x��3<o��&�,sΤ.q~׼�P3\V��39*LZ+6U
���F�#u��w8"�����|&?N�^����o�x�'��ŭ�cQ?��3n�7�˒du/^���P[k*����jO�>uv�j��/"�K�{:|������d(��/�܇�+{^l���v��1l^@�D��՞�ͨ�"�k���;�1�V\�[y�t7����MY\p�{Y؈�=�/��F�pT�����kr�CG����S�ړ\鉻υ��X���?fW��幓D�G̙�<�@*�ߵ8ݼo3� &���W�8:5~�����&��Z��̵;��� I0q�CD����X�*`�F����:�Cߦ��WOÁ|6�+ܱ$���8*4>)�]�&X;Y^4|<aN8�@*E��YVϑM���� ?~&��+��sU(.6_��Y�]���ƅ#�j �c&ʖ-kW���I�������X�X9�G�n�q|��P��c	����V�ΰ*5���$̳à��aܧw����&}_�|�`�]g�>�~J�q(|�1K���Y� �<F!dA�r�y�w�G��㽸��rѪ8T���B�f��[KX�I�3��R?�̳��Ɂ��H��W/*���6<!k�>m�|��E��T���3<b[ҢL�
٣��:˟�r�ݨ4:��:oۦ�±z��LI�疣��L7Lk�깊gn����ŠQ���'6>sp�40��^!���PQ�'ľ<鿱Ĭ����@�S/�����3��[0-�QC�X��������^�'L�"ֺ�mN�"�O�O	\Q����LR�լ�M#hti�YR*ؘd%��X�9��eع́��Q,�jT����X�4o���yr�S�}���M�
��CƖ|�r�����c���j}��;�n(�{���4��9�UƿU�N�4��Or|^��UVg$ ��o׽�Fj6w�s!55����;iR�/A�ͮ�O�ǝ,��9vf"���]��ħ\�[���Mj3�U#I��	G[!�9�Y'���Gd��=VV2[�0qbIj^�ua�B��P�]�������N��)^'�I��g��	@jv�h�\��dO����YA$��� �2��TG��ZPܾ�2=�B������#B��Z-JgWi�h�5g�����ʑ|�Hmf#߉|�ڻ<�m;2N�|�"��Oq���IE_���jc��R���$�fƎ�.-]�w}�8�ƅh�.��~"T�O�.q�'~ k����p�*��MZb��b9�͊7�v�]}�����,��	�|jSFT�͓�v�n	Ni�$��Sw`���2�d� )}�H��Zw�@��~x!�Y��Ȥ�����?Uf����K�1��".-���B������d����� �Y��"�<	�t��sQ`G6o�)[�$:��Al��(�GI�+�nz�'�	*[a12}x���wz�\�n��>��/����F'��J��O] =�{[{���A9M1�P�LO�U:T��A��tAg�s
sX�0yqˀ�,��0�^���m�=dƒ�B���	7+V������O����t�Q����~��G�T��W0D��)�d%Y�Y-�v�s�������Go�`B,M)�Y����W�]G�n.���k�$���(�
X�m���uTP�
�ac+ ���d�b�8s��fU���X.wC���3m}�L>eB6�$�EP�ü��f��aݍkV�y����ض45�i�D�
��;�6-���
�"+��F��Zf�ε/=P�V[<J���=a�ν!��W��*w�WP�?MY6M��2�j��2�I�bR��� �0�=�6����	���
g�����[f>��uHh@����$"��_v|�����? �I+����I��~�>�o�3�4l�_6����N*�:������X�B��fk��r'~�-ȅ��`����4��]hs���jb����oŭ��$�Γ/��Sir!�u����ˤqh��ڢ��kc��Hޅ����a���*�iy>W.�����T؊��R9c������=��ߵv���n8u,~3��=f���}~�\v�P�5�5^W
�#�IX�l���N�����x8��$���"��Һk5�k�aDH�'��i�����OOi�!B/?,sUiբ'�1�ׄ0�6�3����SH{gb��t3���٤��l(�j��y�����W�5�Ŧ��Z��HwJ|a�b� �7�LR����~�7��iflY��5�]��͈⇬�pm��sG�N&q'��.p@�T8H�.���|�ef�q���f����hqZ��Ut,V�]�xK����0x5�3l@����"�=�c��u��^B\V(x�GD��\���s��rt�����ī�QRJ�����/�k�x��j��T�cG��l�=o�L��۞\7���)lst}���%���P��=��s}$a���$d�!-b�қ� �R�	P��X��A�@;��ںe��I��9���;a��;�W�xCH�Anh^�c�����ls{N�5�[-�_T`������G��i�ʘ����6M���ˁ��q�?{X=� ����Ʀ.�9Dm�HrU��϶�-I��}��F�U���d���O��`�U�V����B2X�`Bc��i�	(��$�������k��k����eyQn�x>�.��X�}�@�U!�ˈ��|'��\A�:<W�eϚ�cO��2-�줿��g�mƃ���k�b��r�J1��S�s)v50�Kd�)��H��.��w�v��fW!�a�8��z�8��׆L�b���1Lt��4�fH�⇂���x�A^4��T7����&E�+YXA�� 5�i���Z�Ըn���+��s��� !�j�5:�ck8��F�6
��f]�O� ڀsR�
���|�3M"����5��[���3�"Кj�5�CH�U�������v��Cs^�,xW����Ϟ.AQ��zW���@Y�^�cP
��a�4�փހ��6��(�=n�9 	��P�iB0b�Ū���z�a tDt
�^����w3��p��	�o��� ��~�94!��B��
~��E�WO��-h�v!�&s�	_Q(=�i�G����H�3��Ɛ�J�H},���|�z;}t�!45[vwX�.�� ���!@�N�e�-�~Fq0�6=���S�H�o����_N~v�ަY��\<�W�.����6:}%���C\ֲ=�Z�rA\ lb�{{�� w���w�L����v��Yl<Ch
�ޞ���C>z�Q��+����g�7`��_uʪ��eY��}F�͏W<y���-������I0�P� �jh��6�=@p��h��_�N��@!a���3k���Y��qCV�G�f.}̌���r��H�8YS'�ޡ$�J�ܬǹh"zL���g�����3��ග�Bd��$8Wʄ�~[��S9��6U\��ha�\��I2l�p�E�Pym��j���#��d�o�fg��w1Z|��L���岸��}ZA"�O��h��@��M`���f�?`�#�#Wn�U&�/���4h�g��u����(����>z�{��H��s3_�ף��S7˜R+�@
�k���\FW���#��Vy�E^l��
3���'#�Q5X�����q\Q��&�(���=����� ʥ�&�`���4I�屆�c
���:��=��^���o��邹9��Q��G�*R3�gqOj_!�#C���o���#���=����I4�`��Xx�R=[gz�)�;�g�+�[=!��xs��0q�M��W����x�񝶶:�~�P�N������l����2�����f!�����U��v�Tg㊱��{s%d3w�ec�W�ܩx��MI���;���!�|�F�B�y��|gG��zP�pn
K`����	�{&s����{Wk��opi����4Z����4���+l��ҟl�~@6/f�[��ӳ�h��kH����H����8aKt�R��J=e����7kV��(��vH20x��{��0�L��b`~���&Lң(q'˿�� ����	A�+u�+��6����]#N`�c�_�ů��mQ�R�GÆ��
<�	�!&F����4��m���쳝'��ߐ0��Oj������x̰f�f�t2'a�
Mb�6�CCݏ�ƽ��8c)\`��,�I//V6���������m�����в�q���I!=+�*4R��}�1���Pm�R�oI����9��5�p�}m+��d�4=�4���&ꎡ���g(��g}�8"�&��_���jAo1�4^q	 ��ڂ�U��b.��.O�p f��{��O��ʫ�s���V���Z����|�=��AN~�z;���u�T���q�`��:Kb�0�R#&��R�{����`�Ic�j���8�������)��u3{|[�ݦ����n	���Ox��̓�5k&������ 8)o0 l�F�J�>�C.P�0��C����;t�P�<������ʑLd͡l���+#ӂģhH,�Z(5��ɳ� �i�8�b�i>�W��f���a��c@��f�կV��ғ����1n��b�'�m�b�P��H����g��@.��Ze}��H�#9w���|�`��b@�=+��2+��M�rq�1t�yE0sh��(�Ƭ��"� ��:��l�9�8��C����ӿ���z�r��&D�ξ�A����41 �����A�^�kA�=\/�"0�3g�a�R*�]3��Ն��[s��k����\L��Ռ�;雅�ʞ��8C(��!�d�Z-#"�"��x��o�����~������-������,�s���\��c��,	��tj��<���̙ �HʼDj�yћ$K�������!�P<'�[�,�)���
X�T�,ke���G���M'�T�줯�n����*��ϡϲ��sФLa�O>�޴FJ0@^#�!��z2�]��E��Z ��F����M��?2<4U�������.9K֪�+C��#�/8��2{EՒ6�Do�<TgF9"b$Ou�7��a�Á|'�t���v�ݙ�v���LI }�Q��hP%7PEaW}@��^P;Al?�W5����E�ԡb�2�ԶD�y����~�?�����kn��c�&��0�a�3�r����1�ܻe�&�:v��~D4*�p���=�֫o�v+k ��꾏g��D�S�W]�$pg#�ڥ��6@�����K���1*���4W:�P�.�7J�����}�<�,�b@ng�}�����84���g�gW��e��Wꦉ�ґ2�My�2ٽf��$y�'筸��*qԪ�b�)Dl�@�@)���C��K�/]�����v8�z�/	�v��I�x%���m^���71ɹ�EQ��������k��3Ũ��-e���|�և�#ܘ[��-%)��� 9�
=K��T(�����+�M�K_aѤ�R�oV�/�'sb��
ɝ��j�|�О�"A����"��dAI�O��>=[O��������J*�$�A� G�B����Χn�G
ԉ@7��v7��i��&�������^���{�[�+]���S�p�V|ۄ�+�M���VGx����i]�{�u�j����d����J���y1�k�0�����=d�茟]��wMSA᪻�d�[.�3*|!˯�t��WZ���T0,'�.��"ϋAPj+�2B��Wid�2�_h�[&&�/.�HD� �:-;L���N�J�^3)��k�.Z��X�jb �%��bG���u��/����e�*7D�h�r>r��E�
@Pw�Pfq�y&����TK�����s�ʃ�1A��~���VJ��Ď?�v\j��P�Y����f�Ǟ�\����S}��+q�ѫ=l�-Q+�#�$��D�W�1�lk��K7G ��Ʒ�#ޡgv��$�>�(-χbh�H,F܋*f��5�����IQ���T���F�3]����m���&����Jk��Sj��쟿J�3������v�ϊia��R�n�z��vƖR�]��"��~$��0�8:ߠ�8PU�r���K6x�WW����sb��<ؚ%��[�Ĥ.#R�,m�O�.�����^:����!�݀X5�nw�AI�
k��e�=LQ��@��A��;�]�7Z "k?�l�(׊��`�9+B<�
�^f,����n��\������D�tz��L'���X�.��n�Q�_v&NZ�e�"��Lw���lrOJt
�Y���:��LE_�R��hZO �a��/	)z����*R�u�A����|O$�>������*(xo�T�GL	�U������vI��܀Y�Q��V	�7:��3�C�����.�d���_r����%�hH�h���֣Lݪ�*� �sV��$\��{�<\��k
kZ5��U2�<.�u">�~7,� =�[�gX���MO���M��&���_~s}����pNe�"7�O��"��
�l}ɷ>!����:�L����d��={��M#ծ��
ѫ�Ot"�a��DΒ��u������g���YD�z��o����F!���
#t7����%`���o#���N��u����:���1�O����H�����\���G�_�)k�ċz�����铫�g@
�9�do	_K
���{���
m���^�Ea^�\;8��6�`���i̹��W�䀄�� Ff��L�ư����(=�#�R�%�ԙ����o0Q������^���|vJhm�r@MUݩø��ڈ��G�z��/N�Q.��꾔����xi���.Yx#:v�ʒ�,�r��Ymϋ`��;���$�������[$Q^'�%Q��|��6ʯZ�@^ZNg��J̦�������f!� �`�\V;>Sή�K�{@I�^6�a�"�P�@�����P ��2�y��s��������HR�ǽ��;9��s���7�!��ݟ)�>�}�0�Cv��`+�p2��w0?&>��9���)�����_�e�J� �5u����g���$s|�Ε�j�b���$����9+q�:K2דS5$W��VՋ<'���:f�(����TEyT�oI!�	:�!Ɠ<r!Zq^��2�p������*�4��b�ζs1��KD{����#Ks��H���|�!;�<����9>����?���9���CzR��H�+>]��ZX������z�G��e
�ⳤ���9��6�#x�+��}�	�mɋ!�]�hs���.��{5AKm��沍����N�G&R���2���T�1���)�n��G��1Ru <E��e��%<�^��8�Q��_�N�V;JY��A��[�BC����$���u�����Z�?`a���_��CC��>f�1�q'�Q}���#K�I����ɕE��tu��`��v}�.v'�OC)TJ� l�� aD��l����O��c���+؜A�Rz�Fe���!K�8<ds�A�£>%�Ņ�����YBH���^ɠ�'K:1�S+�� zU��6D�M���vܖ�v
�ټw�hd2o�WJ:�cxk��M8�� V��k���5a���l��{/ e&��^"I�(����-zӳv=�p+NpT ��I:n%|'�q�.!�����U�tG��������b�oȞ���u��6����t�����W��o�	�Pd��̚��5�NYk�6���{�g�n&
Z#JدQ���`.�[A��dL>Y���KW�8Zv�yEM�`>E��<�2�Q�YJDɺ0�C�
��qޗ����/��ל��?�{�<�]CN���Hܰ�_[�:�H��Y�+�\�Y�n��>E|�@�؋ �RU_���4�Τ��1D�����י��3�6��v�����.�Y<߫?����k�FNy�jn.�,#�ىIR�"�Iyw�/�ax��UlձZ0G
��^����P�<E{`�_X+�4?���w2xKs��+�|�K�������}�;���m�^�@*��dJ�IO��i\���ULN��	��e��+������½u�(#��j1�"�l=ܐ��NK�����7� 
���c������\nx���]V�樧��i��7��`=��6Ux���\M���k�������;��W���pW-)>W&\��R�-k0E�:d�yWM�f�I����kL�t�;� ���Mj]���/�����[��M^�@'T�f�l((���¤Ӭ7u��]��v��
�7Ql���h�s_V2�1{�*U�/����5Q�D�D�Z��A��[�?F��	���_kO��g��Գ_jh̛n5@�l�����>�׊���xi:w"��>}Tj�e�(�+'���AD/'ZBقg&2]��- ��3�#��J�Dُ��ODy'|y�"c(?�}Rg�� .,\�l�}>��A��LYaD7+[��]V�-����2�.d	zѡF	�Z��5�ӓ&�V��#+�R�풛c����s��U���YF��X�L�>���U�V��Լ�
�Ml��T��JNŝ���|�d�`��k��#�L����z��.T�'y���{ lÏ��!�|_g:DP��i�鮥n>Ɓ���篨7���d�BC�z���8�Muk�WU�ऎ��o��cE����8^�;��ׇ��i��<���C*�;5���Kd>��z{�D~֧�ob�x�MNR���0�9��"���/�$TލR�p�ʮ0`�:��)�{K���ԯ�����@yq���!���E�e:oJ��Yr1sj��;��a���}��,���kz�?'�x���\M�=�|3��G���`�W�es�I���j��� ��2����!�}pF.o>k�z?˸l˄J����d�	��F��8� A���!�����w/i)Ӥ(�����l7f{�K�n�*�tu�$�J^��k���I���ܜ�i�������P$7�c;n�Q@�;5�ڪ��'�>Nߋ'��4����x�g݋W���{�%���I_������C�#�
H��Htua-$���I�4H7dL7˼�� \c���KF�?����"ʪ�ar��>������#�=p$��E���"��Dd+���ʠkDD5���|���0dǡ�P�C!��V�)��75-N��r�1|G��{�V��AH��t�y���eaۗ��כȕ*Sx���+�y���b��A��g�uXg�x-8N=�B�淪��h��9	sC�(�,?�	E���{�78H��}{�^.=��[�����l�<b��xR����6���UMD]ǟ� 9B��`<�l$.�;�q�`�~���1����χ�Hiݖ���ߠ��<l���|�m0�i�m_��9L�̪���*|�P��QZ�&޷!�6�'k����P�;7�P��P����(��̏A�C��I��Fh���pu��j�9���� �<�jGY�Ƕ@Ndj�q��m��1�|}��񋾿���O�� ���o<HPt"�� ��a��q�=S����7LT�]�u����\��_%�B�k��&a��G��:������A�O�	O�?���:F�U�5̒z��G���68�N�Wz�h�q���*Ӽew	��������v᜸���U�a�Ǯ�ݰ������K�jέ�H!�^�8�7�Fܾ�a��������r��?�x�Ο��C���������b���T�=�I���{Eu��]l?-..b�7��b�Ic2y q���[y��TdpE��j~��Ef.��T/ti5��7`.V,��n�@�6���K`2�]=l��n��OLKf�����kG�"?wv����z����{/PH���մ>i0��;<�<Ơ/y�e�y���r�q��[�������de��j�����ɻ	6 i�l[|U	����J��S�t�A��%�����#���>}�4��ke :E1BQ�JVP���Ȣ��#ܢ�d�����bi�8���g��U����0b�'�B��
�E�SY��`*f��q���Lm�L�6��<C ���V��\�N�MY�9@}�}����~JD ���0+ůnOH��0�ĺ7/E�k���f�mF�!�IqD,[ ^��&t��Ʃ�\��Um��Տ.ԄL�xϘ9L����b��s���~L=�a�dB������&��4g�
f'�(N*4Φ����S
��Ê�d<���"ͯ���ݻ��;���g��,h�;L����8�:�K��v�ɻZ�)��4���I_DW2y�}qW��������?sJV:�����3�P����+�m��Yd8�&k��֙�&�7'�3n'��"n�}�T�����C�}�s	��rE8�����2*q������
L�w�-��،wM |Y��[U" �eaosȔ�Yv�������#���l\ [?cRk�|]��4?d�aغ)�_��q�H�I������Z�A�B�G?[}��@��P��=�O�&f��5�Ad)�jetE�y�tt�ԝY�令�+6�L�fu6i�
2������F�ݟ1	�\@%�|Ț��%�D�04����tIQ1C`��\$�PH�Y��-��a���D?��f^�u��j �eW8S>��5��O��[8ُ�Ua/�oO8�/pI��.�`�n���I�^m���^B<!7F�t�Q��W����}��6�XM{$l�F)�?2�ڍjě����6��I
������F��[Y�*���֋�j>�N���3i	Ff6ĵ�!Q���KQ������D�1  �OtC���&��%���v�#qT���\��fTe�����2���IM<��0֭F��؏�89�2�j6���	���B�4&SnTK�t�;v���r��v�dY��q�;a�)��O~E�^ګ�F���wwX�@/:�	E���f�������An����H�������e�R� +�$݈r����� �p0���13VcG��������h���%2����dӥ��7�C��C;Xh���X$�&���Nκܩ؅��Ŀ���p��% ��2Dm�g��4P� Г<���N�D-b�yt����R*ʫ��ձ��� �[`�Y@We������5�J��M0u�g��i�V��}�`�[d�I�gA�L���:Xxp�<aP�G�f:�=��������R�@��(�/$����^���E����V��OB ~��v��pu9�<�ɔXxT���L�=-��N�.&,{)$yi�.J�H�����<w�#��AIk�[�7�tGvSM�t��6��0ye�rN���;g6���X�証�����1�" ��U��}v�;�fwMz�nΟ���O�|i��NSO�%�]A�i/<���e��ŅB��4!u%���[*^�,�ky��Kq����4���k!myL����OQ���9�/����lZs�W��^��3��4�ް�5��?����Al�U�ҁ0Uz�/�^sO~��y[5iz��+�6����h�1&���c�j���_5mVq?P�S_P���=�� �c(^zP�kD3�|�}���O5�Mpb�l+�v9i�L�1�3[��T��5�H��:�i�f:�s���t�ǥ}�����i!-�t'i=�)I)(x���D�9s�5�͍��o����v�pn�3x�1����6��,��^f�a��ey���)��������n�6�����Fw����;&�؂�cz�̿g�����`%�B�QG�P9
=�_vԲ��"o��Պ��L�t5�|Am�l9�!e]��m��) E��U���i�����+A;@{���Gj�#ub�s�_��3��g~+�d��Ŗ�E��\vT<�Ɵ���Z��B\ l�3TC�����Y 7���,�^��Hpv:W�Ch����a�$(�ǡޞ��RO�6�89!��Ї���w�Y�\��\1�zl�`t?i�	�I�%׀3�vNݝfX���Q9�X.�@C���Ʒvu�>��,��E�>;�/2�
QMLf�9�Q��ӥ"�aį�Y�7�v|6*D��-�'�x#�Ψ�JǇ.H�4t�����߄�����tl��q�0�+2GZ҇y˵f	Szc��p��e�7H�c���q��l�[���(�N�����sq	V%�������ҵ���u��iU����Q;���^�	h�RVDlHiZ<;�gO��2!3|��&}�n{��>���S�-` &�XS�U�����qՠx��8K��urG�'�Aȣ�i
R�z&Ԧ���mh�&Z�써E�ab$r��b,��Ū*���3��,�*m��>*y����z����A��sK��3m���^��2 �a�l
������M�i�dF��X�����1�VY	�>�9�C�b��牚�I�Jf{ŮiՖv7綤���U.���Ǿ���;
S�߽[���1c�n����%�}��r Ѳ�,�����ݝSVS��c5�N�5�h���0~D{�O�㯴�Zz���q��1�cۃw��Q�z76��BZ*���$����Ҧ�q���B����m4�64���v��%��F:��w#%�q����t��>���~x���L��k�|G_�^��~��&cWs�_�#�ݽ�mQN@y�,�/^��O��˯�n��l^%>�ĳ(4JcC�c��!�zߩ���U�;�sH����_S��[�X��q���Q�i�f�;/�T"\߳ܚ�=�Y'A�D��Sj��4��*ǽ�;��ԽK��}Gw�ׁ�S֘b����BZ`��g��.;9kz{�i�>������� o�o�Z����k&M���oֺ��H�����m{�Վ�Ѹ�ub�O�Y_H{/lW��g�bZ��V0SX́pF�Ƹt����E`��?����U2�5�Va�����iUF��G�C��[��sr@:F��a�����s)��V|e�,d��%	���P�f�17��)�����t(:(����f���c%��������F1��L�C�5^)�;��t��br踴,�j� �9w]��~@�jQ����
�\6�ڞ��ة�X"�����Ǘ�|хO�5���_wo�D��_>T+Nz�2T�Md�s���W�7"��
�'���Jm�u��z�>���L�\��5|�f��ⱏiyޱ}��Z�L��jօV��Z�B�se5���Ͻ�~,��n6rY���u ��D�"R�]��=�J��4hW���qv��4��g��xӪ�2�O Ə"^�,��ʕ�zǔ����j�vm������M���j�fp3Hз��"��7���3Y��.�@&<[���#gҧS���r�x�!#hrv@�y"a��C�@���
�������8'�zn�f�@.��=�9�.Iw�61\��m$EP��=@5Td/
x�8���̔��`��y��hn�:;�2.�����;7`��b�WL�62�(�� P�&Y�?az�Q&�*�:�D�$%����!ʸ1>9K�{�^����Q��uL���k�����qC7+
�������X�`S��9))�5�R���Cɏ��vح���<�7�Z�����1��+Qu��x΀ �
����2{9��a��F#{}6:d�@,$�ٷe����Y��i�<�#
��#E�~q����s�DBp����d�j�q�wc.��Y6+�L�{�)�y�v�<R�F�⧙/}5���S�{�kL���A%z�Ybd���~�P	���ƽ��!���hq��d����L$�/��^���R��͟�~�@�q����/ӊ�R�K��Ţ�̌��Vz�ं�w+'�Ҏ��gs�����R�մI}�Ts�
�R-�&��Ht��y/8]n�߉��P�ik^�׷�-!�'���ƞ��#ڦ
�K��o��?@�D
���g��W�U4*2��M�1F!��?�E�\lC\���v�A�9�f=�P1��d�sՑ������<��]A�'$������(\F��?3�A�.s�9.����鼎/�E��6�<�l\'��E��*�����H��3b�Ď�j��@u@���X��W��Cʙ�>6k�@%�#*��LJa7�[DV�ٗ�Sr���JQ��6O�Mk~��-��[�Z{*��>��#g���Bn�4�t���EU���TQ)���b�7���l,9�5��4
�?Q��B0����bu���^�5_����)��n��C�x��-yPEZ�9�~�>^��}��`Ŵ����K�<ܻ��Pב�dL)��]�K>�l-\��u��D�:��O�_\J�B����[�CS��Jw�?�E��"��O*��8�'0*U)�_8�:�&��è2�!��O�Nه��R��8o��p��D��h����VVv�cv�⫷���`x�(l\���uDF!4	�����
�@��f
o>�):�
se�`~���Uafm�7�����aO:K�}~?�`ᷳ�g�򺕂^�C��x ԡ���R��kĚ�)x��J{�E�6/�!+�.5Ϩ�{_|3LW{}/K�-q�o �T* �;A����s�$+������ksB�I�{��K&Q|S��]�e�[����w��NʑYb{->H�|�4X����֮��J�`"O$x(/yH@���ڰ������Q�S8�7�`��~��+2�����6�%8Ml�	�i:�ٱ�9���@m!�d�T�'���$#v�}�m�"�A����A�gБ)X�.b �06Q��ӹ����ׅE<@�����g!��'*4~<e��r�� �8��?N��:�F?K��v��I�o�~��.�y�^��A,�m)NM�M{ �KS��99����E���U��J�ߝ������X `�z���{���D��d��j��:���&,ۿ0�<ﮫ�j���#\������=7H�3U0�*-���VW�Q�%G�Y���H^%[�Y�=��xU�M�%��S��B"�#㜎�C���^�k��+?�QO�B���]9֕%��-P�x��×k�����L��� 4�����[���'���orH��WW���a�R��M������4j3-������Ǎ	�/{�e�w����s��^�\�٪�7�v���\��~�g��c~�YTb���eQ���+.�*�H��ښ��^�����Z����8|~�Y��M��4���O�fc���'�����G,n�V�D3xe��V�*5�T	���r)�z�����>qx*`��}�9#���ip�y�՞��$(`	Zc��o�F����ot�����W6�hV��C�ZA>�<�ÖQ�Why�1\n.�k/+��M@	�Ǽ,��`�l�Ny�^D��,���F�Fo���A�3�T�`_j=�����!�1G�����#���sx�w���~8*�?�MH���V�,���i� 2	��7�Ҭtt�7&<����p:ɯ���/"V��w�o�!� �5� ���6v4�}2[5�Od����.!�.��86��j�V�p~�z�6��eb�gdk�5v�v&р�@t)�Z�X������*t���9�WD��|7"����c_B�FR����
"`yx}���� ��i�ӫ!��~M�~����~��86"1P�es~�$��,<�=�(6�i��"e9�θ_���]�a���c���p��?�!���z���۸���K}�_ޕ2�s_��{����w��l�k��6t/���26�$��ln�K9	R7���^��gk�����	bJ��D�sni��ǧ��p�=ٲ������A`��V���bv4���ǀU��)y����R�b���4@������O����?�>]o�_bj79Z"xj����(��y��J��$;��SmWX�'�c0Y�؋}�I{C8R��}y�����f�T�T��(�!����<�@���N����/0ՙ	M����&�&�m6�������h<3}i*�Ũ�LU�[�w���yzMZ\-ӝBD���`3<Wݔʔ�N <�\c��Е�M�B�Ge7;�L���r��j�`/cj����1:|1C��\�`0�d���$��C���p��'o�����(=�=7b_ <��f�"���ph���E`�K���z�*�	�*�A�,�������gV=�|u��l������?Ȝ� 0���v���A�&ρ�
�7��	Үd�и�~gj�5���������:tدJL<o��t�U�W����q�g����:c=I��s���[��̢�&i5��!��+�d1	����<�X�qd�m=�r#TKF�6���~x��o�P1��hrj6<���+��h�]��(�n����҆�-=�q,�s{��_���!1E�7����4�oH�
�J�� Y9���!�l�xd���st����0�XlJ��m����]�i��f���]�xv|�%&Ves�*$�߅�_$M]�;�:�{UK�E�t�t{����~��:��i3;C�O ����A7�V�꼌��8�F�1��"�*�@�<~R�72�����K��J˨��H� X]�)���W��}q�W�Ŷ�9Rh*�&�؎`-~_�6����{��]��
ɭ3J�W��q�V�wk��݄��#��b�:�7hَ����2Ѧ��b�V!r.s���eX����$^���ȑ����8P���i��{I~�t�Z��:����4���"��29~^�v�2@d#B8kS7\i����S[ 3���ew��^��$3Z�.+��{���O5���,1������F����Cfq~�U�|J��V,л�4�=d���5%��}�[x$��J� ���U�S��I���XJ�ԑ���IS����/�Q^v���`E�;f�܋��4�W�1��-=4�L�;Pܻ�[��h���*dL��E��֭ ���;�����P�ƛ��c	w#
���#n#��{���v>�@vbL �~���[���؞Ҭ�O*�<o=�UWr�!�����n��~���F��uum%�i����$���&����:�@n��eY=���-�OeTV�O�Ǿ���d�h��b��e����H٧�bYeB�^$b�h�#��ǋb��
+<� >�N�<�zthj��Bj��������xw��t{�tl�a����x �Q�:����m����B�ڝ?��d.�2v�����e5O�)We�_X��ť�v9˲?�2`+>t�in�%�nH��0�J���*�D�Cx�7n�=ĩlK��!,�"�
��3b��H�f�`hʤ��|g����zJ�y�BQ���P��0�#�[.=��b���+���a�E�Oߙ`G�$�7��"��!�-����n���;��Ik�t5�C����t��q�\�m�7��a��ci�Mgh��9#~�O�����%�F$f��[����o����D��M_ib 5#�_*�`�Q�	
����ha��+�'3����"r�m��,/� W�d��e��WlM�j�@5`���Ta�2g�췓���]

5=Gz[�COT*�+bV`C�ś�$ۺ	s��$ز��=��U}j�w}B�4U�qm�s��J֍@i��:P]�5!~�N��0V��n���Z����m��u'C����S�������٪�u�=w�4�\k^J<�,=�b�$S����fTY!�4���?��@b|�6JySd�r���v#�V�f� ��"A��u&#/��͓t0?�dz����b�e����wv�E�Jk�?�������D�X�X�J����GH��2�ެg�s:ySW�1C����Ӹ�'ݛ�/М��U�؇��%�p�g��L�`m=������wx������M�#�
o���F���WygX�̽�E�:��b���4s�,G�K~L�������z|���j����Z��R�9~#������/��J�+��p��(�L�|�����j��R���̗Z$���8��$g�O�φۛb���<:�K-��y��_�-#���O�3 _ ��h��k�_�x���e�'	</�/�d��r�s��[�8u�}ې�)J���P˪-�0+(���%�����������s,{��`�7#�݌���L�n�lv�(R�Q���a��V��'�:����o��Ѳ��-կ��������ڲǿ������Z�D���EPwshtY����O������w�������&�@��V%�i�J��vY{~��}Z���?��4���! #��7]Pu�eYg���U�?�=_Y�C�A�]ݻ_����}�5䗑@`t)a<tW��Rq�)
�.`MH����?����z :��[���� �L ���֏�����	���/��-Jvk�$9��Sr	Pr���ڂƆW�u�"��H� �ϡ{�&/�z*��D�n��wA��*��cpf'F�̪e�����Knǥ�R��:<#�a��0#�eOD7`��MunQ�l^�%}[Q��>�|s]W�����b���:��̛W���N�����U�����Mu6Ac<�d�L��p��FR��lt:N�4.�mA���ۤ9�w��3!_�*pc۩�i�ƒf�����s<��n%QZ�-�Hk�h�"ͪ��W��-��J�n�
�3�:��ңH����h�?D��c%61�i/ب)9�;�IaL�
�H�4���z���ùZF�c���������l���te-��jO��a��SQ2����)�hj@d�+���s��i(}��h6�=��u��~�CHX���TCO�]<�>�����1q�|1���R�j�������Ժ�x�w�ĩ5,��J��iΚL�̑"S�u&@�f��7l.��
q�8s��N�_ a�|@����q|I�~9�a��
lɮ\�>W_�6j����� ���M�ԕ5�>D�&��G7��Z���7��Koy~c�s/���|�m6u���]p`a�vZ�D&"^�!A��9��wY>��H2]��01�{�\ؑ,��uBOX2��|A��Ǫ������
���=b2Eإ����%I�8D��D�~��6���5��_\�,B1�4Q���&��/v���(�:cO9L�8I�r�Xp�>�U촸M���Rg$,[j�k�[��m;9�J��=�ɔ�}7�i�%s����A��l*k�`��h���w�?��ki,�Sva)�,:L
9������1���U�M�Q�A�b�Ӏ]F�)|���`��	��$}E���Q��[��(=~S΋�;1��s�U���7;�y�x#�`	#*�X#Ad�k='��9����)Jq4����Wcg���1a��vߧ�ߕD�է���?�K0�fq��~�s5�($]STÇB�5Q�m����.�aF����.2o,���0��s��G���2���a�(>Muo����RNjK�m}�h"C�=�W5������u�ZK��{"�4x����@U�d�+� b��Y��_��ʪh��1�q�h���k�����I-�	1~�YE�[�p�A�`J�4��F�R~��Ñlܠ.H�#�s�W�.^(c��&N("8*2��9����{�#�2�ql�����3g�����x���1����v[{�%��[�� ?��sX�p������.U��*�u���xP\?J.�+hH�U%=��TL�ǉ���FB�<��gC���o�Wr17���m*��u^l�ԝ�J3!�rc��ԕL6�A��=~h�gP��2�iG�d��XX|u���y2��;��4"��!�aRʲ]���~?u���۫��g�8{�'['�YvB9�à{J�!(<X��9���Sߊ0�Ֆ��	���N���qv�e(��~�E�_��8^^M�An��p����Z� ���o�|���Oc�Fa����������L��C5��0Y��)��	���wt+Ŭ���'�Є�������������(��aU�,��o�ӱ{~��tfO�&�/�Lͅ�O�Z-|�]�b�I��Yq&�ǚ�#�ƏB�|�������<�Q�7[�f��Uq�x	v�w�nr�#�Ӥ���^�1�G���%i���� �]��a�T���ŞB.|X$��\�
0��#�Z���0QŨh\����k̕����e��y�p~/����ڙA}~���*#;��.2�qz�j�o��3!KN��}p�֊6���z�����T�Gr#9�OKErKcg����&HN\���[�,+�AW��i����i�h����²�F�z�ɐ�$�'����Z:|����2����b]dg+�؂�H2D�������̬w*p_�n�@��Ӫ�?�`NZ�za\Զ6���hF��6��	���mk���y�C�t��Tt�=s��T�#�`�fͤh=��!g7v*�.�� ����|�h����g�����1]]�	C���� F���J�8)T��PG�a^��Rq����;�wӲ�Zm?jq�ik��e�������"s���-2�]���y��L�i4S���?Y
�@�[��&�	w��< F��"���7Z����2խA,�o�����*"��(L�f=���/lL�h���%Q\���ǀ��/���V��������)�n�<V��m�V���^���q�./����=���dO�e��Vu!i��|c��Ar����	�ZTm�B˵�z��l�ve߄�Vs�&B�Oh#O���B�& ��g�᡻�"��L����[��,��b��^��� 7<薂����C���b�ڟ�"~��Y�-x���ٹ
�f2�oԬ�ё�J��o�L�>	�z�)�A�\;�4ࢄ��ylq�t�-|��_�a��($���JE\��_�����7)��hH ��{S:G2�O�� �;A0��|Ɋ��@j�|�Q
�E��R��<���jkc��6^\hc��x��a�F�D�}���d���"��(��] �j���/��\T
Xg���(���{~a?�e�Z����:���˖	^���	ꌬ�;.��w�C?�^J���� `�ˣ������Y;rU��؞�穐3��1M�QW�/<�i���Ǣ��m�ֶ)Pc�>�� 3��ӠxI,Յ��k��pj�LmB��i��N�n���	]��i�C�\T���㸤{īXw�n�zOHS�X>��1J�A�.�k�P�%`��6@�)"�x��r�2|�e�����Ԛ�c� {�B��sCSͶ�;��`��w��y�!�Y����2FwA���Ug��ޱ�~l"�J)����q�{��U�>���&R��e;�2���]ȼ��	�	�N�5OジH�}0K�s5�6�J��
��b�&ʆ_AEJ��)~�3E��-V�x��y�C�l�����c��f+β<K]߃��9�_1����K9D�Н�t�_�	dzk�L:l"F������C]����M���2�'�p���?��z�k����ɒ�</�P�.W]�R}x�7L;��]�â'ׂ�+c
�)f��S�7�;L�#��� -�+���tr+mM7nh�Q�sxД�h��&7��We��G�}�8��|w�����-R���T��'�ye㻛��׹������k1T5����O0X����Ƌ{d"����%�0J8�OX�9rKS�TC�M�wp��u�{�*v��x�S�3��,e0`��ί?��.U/1�,�@�I4��2/���I%ޅԾ0pQ/�(���5�C H�*&y[?-u&�$u����Ѩ�NXH
Ih�'9�nO�b!S��e�.͋��}���\
�f6<��O>~�">UHK"�>��>��lX��4�jb��l��MD�bW�I{�]H�������]�ߦū�`��PRjv��lO#&*փ��u�\�Q�^���r2��I�io�K*��ca��"<�D�8�3�^Δ�_i�"k�t��K�P���>�*�+�o8�;I�B��
:h�|W�~�3�rjT���-�!��o��L(l�7dV%G
��hG�PE�i�R�AX��S��[#�ni��k����7�2`Y2����ik�F:�5`Z��:(h�q�"7F��
0�2[�هH>43�����Ę�Vfo����!���%H5���`."
�����0#�ux�Z��W<^��s`�,�`%���"�.6VC��Ļ�"����q$��!1����;��	h�Û��f@�#�����g�,�a\Z�c�@[��L�s��c&��,7�]�b��)���/��H��D������z�^X�T���,n3��\Z"��N�V��gܣ�D?���8�Qf��)?�߇�5�qE֭�&F�Xm��dY�����ɲ��+�F�Y��9`X6�OA�AG���;�A���%�!��Ð����������7
?
&�6�m�0�%V�Q���z�$�]��I�9�浭���D�!���By��dQ��|@�Mk��zZ�����Cf%u��s[*��Bq,�ڜK��ј�迍��ۍ̨K�ӱA��%��z1m�zO�_��j0�PN��h�4T�T�9��pMv}�[�ƙ���>.�B��j�v����z�_�@��ò�# �M���c'#��Q_7�r���Į� bb�J����������lt�U�&��+�21ֳ�����>>���-D΋��9���Yg��1�Q���{6�����_ ���9�������=q�/�Ƨ�y��n��T�)��D��A���:M��҆��Zp��4�j�*�-�]ܠ�L�(�aȒsfn���"A����h�E�YdE������J�w���wUx��V�����͟һJ��uy����y�¯I�T�(�md������G��e��!8j͈X���&��b�d�|���=��͈�#17��9oM���v�J1w��fUS�yl��>XS�@)����[ܧc��%~���R�e����t�s1*pw�<y����gv�V���j�t(.ޱ�C�V���_�|��u��yʢ�輪��ʯt]@�'&� �I������:��gWh)�L^�`�̔���>s���}BH'I�-=�|�x��$ �:������*�T%�Po������?Vq8N�du���vmȽK��3��A�96s��&o!�/��xƩ�J{���;@(|~���21K-r��E(�y���3�W��+�x�܁��69�fd8B��tQ�i����9P��89�V��va�������ƈ�e�%���=.�L(��2�E.�mFJR3�t4�ԯ��b� ��Fo7O�9�Q���S럙��1 ��1!C|t뎋*D+xԠ�CU��@w�lؤ�\܈�[o���Yќ�6#�<�xH%��#�h$r+Uw6�_�L�@�-���!?#����%��������n,�Z|��̺B0��RYUVe��䂓~W�Qj�J�~�L�ѭ[�����N�l�,\���)/PaO�o�Xk{IO���2�h�%7n<����?J�9���_,��f�����LQ|fd��>q6((= �n,,x�`�6��9c�ɤ�ι�c��b�]��,!���Y���vP�bTtTو�7��9k��G�"
��ZV�]��q�W�e��)6�4J�r�m�5���tq{��~/�I�(J�Љ*��o\x��"��0���r
!��ًz�ڃ�r�e�[j��8��~p�p� O��'�� �[?%�ә���h�]}�K�+9I^z�b����Ӷ��-Ig�=��tp9ee��<����+�CJ��ʟ�.;���r=�#�Ɇ�����h�<c��h�v�i���]�}}=dӂ!:����>�1�Xe��|]e>��)��Mw�=2|?����	Th�^C$�R� �j�!�l�o�����fy��>L+ӎi�,iE��d����o�-�p���!d7�[򀣖M|ϻ��C��t�9����c�+�����!ϙ0��,'A�\���Ȳ��ǒV������;�@��F�rX�AN���qy���� ��4�јu[A�W�|?A%r!*I�� 
��ШKp1=k�:L�B`J� ��h� �w0q����n� b�W��jc�e�Q`�^41�N�"C��B�������$H1�v"[����a���rX�Η�a��ˑ3�V�y�B�Yײ>�H˛e!��a�H�#����qQu	QЙ��t:�^g�5;y�jO`fj�+9ّ�/�"��)�H ��~�\ǃ��Q�U�gNCIoQ��/��G>�]��Y'�r�Ք�E�WW���:G1�a�wh�N"i��N����@Ⴥ|5iJ��K,-��$�X���71��oI+�0WZ���!���l��8@E�f�w����y����d6[��:�Z�U�˹���ބ/�9w��@��f�Fv��M�Cq���l����(�`U���m���/{#�9�G�G)~=��P�0��ep��<�]N�.Qڮ�á	�ݯ��p�����Oe\���Fpjɰ���^����2�9 ��Z+~�,%�$��(�Wg���~Ҍ��Hu	~�!����K�V�	EI���D"��ʰ��էя��h{MUF����匑�A K=\u�P�P�� �M!�ͦ ��;�U MU����o�W�Q�)�B�/ρ��xY˴�4vL�71i'��?
���~N��C�$a|��/F�{��¥�wƾ7����f�u�EXq�s��cqlJ���շ�'�_��2��b_���w;Y���)��	kHs����(n���׾@��n��Mt���:�z��$[�	�I&�W�Vؐ�Li���c�DE��{��Zrq<��&�t۪����Yy���qք&����Z��5#q��J�vA`QH�N
5H��(�C���p���K��������L�$�~�b���$zCpi��N��K���A
�f�t$��V�����mA�U��>B�I�\���x�8���5���b�TΎ�-��W"�3#�fj���6��ޫ��h��Њc��4�a�����s{�D�3��GM���0�)���u���Ȃ0.��Q���6���w�/ˇ���Fc��Ei e�?��ÞeD�B�|�.�
��y�T�aK��@��f٣�� ЋN�+`a��7#��1$$�6*@����.T��u�k皢�Q��`��z��[�}(r:�2[���涮�d�RM^D"�:��>��w��fgu��8]����)ZJ@�$y�;I[��v�4N'��A���o��@��snM�"Q�~�έ�Q���؎�ИnrEϫ��\%|٤�k(޶��	@rK�N�xU�T�K���gNK�3�z���&��;�~�����ʋF�CE8�_7͗��c��e��o�$�~M�y4
�3�Gj�ݪ,�RG?Y]ĵ��W��I�!�=i�����X��|��bEĖ]�a	��H���Ѫ"���M�b�uǼ�`�I�*��sV�QV�]�:d���m�/������?�A%��� }T˥��B��[<[��S;���F�6�Z�.�%S��b"oz?�§�����X���HY��^�����"��#e��K����F�}hP�U|r3ݔ��R�
��B)$(��3BC�.��^W��[��uAf�����(��Ev�2��pJ���1�c�a\�Oqz5C��մv�N&|�F��P��"SGHnt�����X�<�/j���w���׮�ɽd��Y�8�
�n��M)�V��"f�7a�d.�&���]�0�g��q�ݔ��|_KY�#�!���}v!�+�|���p̽\샟�l.��O�G�՛S�Vd�j��U�S�q�����Ez�U��QS����b�RU#�>�N4�b����x,�"�]Y,[|	��Q�@C�z�
י�#�I�O}P��tML�+5�s�W偳�	'�SFmzM_�Z��Oe��Le�Xj�*h�LW��+N�g}xԲC�2�8�P��gNi"������JS(W/�E!?�_zvǑ��qȔ/3���m:u��N�8NR���)R.\�N�$�4�n}���P}�P9�`�N�7\��|�!}(:�j0P3�F^��p�d�Y�bY�˻w�k������d��gAH4p�\������&��8\�*c����٦��y}��_O��;��׏�qv2�I+pX:��3�D�m�Ys�H���Y�e{��#�O�S�Lіے��t�+�m����1�����D�,j���b�<������[���
(�v��U�*�����
s�,r�	%Nق7l¹�cet$^�
Ԁ�&��"�xA�`A��<� �7�+s��)���8��"�[+�j���9U���t���8��ېI������4�+-9���ƽ����n���V2�ʸ6鑑��9��)� ,����pM����H�:�b@]��~����ԭp�s7�>����nMB��=�hՓ�VO�<<�>�5�-��w,�X�mj�`��5[R�/ą6��ߕ��=Q��S<��M��eE(��D/O/M�`:�/�E�z�����*�Q��-���L����t��lmgx����stV��u�-��Bx6ύ:Kvti����@>P2|Y�����U�1����!ǱJ_�c�mQ|=�6�ԚV�bKگ�3��;���i�;��L��'��M�2m�ئz��d.��v7l�n)I�BW7Z8�{W����R��"�T��J�	{��XFX_�J�5��!fQ�C�ЌQ��;H��C��Ў��$e2�-SJ���i~؊�Vz�d��D(��v	�aI�Zɕyx�~�c3~σ�T��Mc]������_,q�?��Y!��?N6�l!t��K��T���E��K�_��̭e߅{m �/C(�����H�����;����2H�q86m#0�->��	A�h��W}�.�V��Q�|�9_㝊Dy^A���[&W���1΁q��?��>�M�_B��K�pu�㵱�̏�۟��dV��F{D�3X�^\
���ب(�����g 5HF����5b�0�����ݸ�2��'�w$����������)ݯ�p+��8���}?�i�����"�/#r�~���(1���D�8���pl������p|c�S�KA�e{�� ����<i�
\.��\����W�S���)0�"N�D�h��t���#�C41m���d�f��!�e����:y�^J�� !�>�Ԍ%�}���SҾA������
M����)�@?�%�ڢ:�{"
���3�>��`Hh	t��w����!l(���Y-Nw��FJZ�����Z�,K��ME	����=ٹ�xҡ�:|b�r=��4� at8��P{�w��2��c���3q���3�`�I�:̈́�h��b�Q��h-��M������$8l�"��(Sm2���n��3����=�
2s�^���V��땏/���~��y<��$�fdf�8�(��{K�Y�x�d������,��-S�<7�V���qM�Ss=f���K��X8�����p�mEp�i���ʥ>�1o4\�KS�Z�zDa.;}B�����W�ȜQ�2(���ۦ�Bu�V���u�.Ri�Rn�\����Te�ٜnb9^��S^ID�M(���kp÷5�I�/�����mQJ{�_�F�4��^T��m�d`��_k�}��C.���X%C��ᚮ��s���8&s�@�xJ����2���`ݍ�?���9�Jt�J�dzKq�D>�oR���U{fB^!���s3> ��"B��jSɷ�{:���Դ��8�N�oǤ�N�,Y0T��o<�M]�C���ݥs���/����(��n�}�������a�~��.*��ezF�+�1=��:#QY<��䨵�;Q#�������kU8f�i�uR�~e�S'ͧ$b̅#J�v�@Bov��s��XO8�T��iqڡ��l���:������w%�Hs� j�&D�]�jI>o��H�+�d0���?����DMW>,�)>�Q�D��0H��	m����]dsqT��CR���)��H�n��:�ʵ��膷,Q���P
tA�<�]xE�_Ѧ|��WCO�g��yg͚�8���eM(ê� �|/F�:�j.Q��]����j`C�S��b:_up��5;`�
�[�S��>&�O�ж&��]@�i�E)}�x�A`>)p�$��Ǯ]����R�ϭw�/cdG��c?]��w��B���\ÆG0���b��`�����j̀�9�2���@XY>�T�^E�Hk�N�^0o�XP�	�:��5N���ۿd��-��s��+��H��c�7��D����j͠���%X zBQ��tE~�[?�!��Q�8+��(�뒟�2��;�7xG+�[ ]�B����7�a�yF���@�/��,2�*��� ׽��A��Q��D�wog�`蕉C6�L�秺��Π���Dè��R�͏�d�I��i��ꉨWO��)�[zɂ�Ќ��ytQ�Q�|A�H�0�y#�|q���-B�t0��{�����
P�[���]�Ѡ�{$�vލA���w/����qL- ��=E-�O���4_�=,E}�a������߻Z� ������}�P�!Be�U���Dv���]n�k����.���'�rO!y��R�G��mr*,�E�r@��i#����I-[`���~�?A�+4�}�M"� X�:��
f����ңt���`ܷ9�B�&���Ϩ�g�����4�	[�b�v4ݤ<`�6A�e�B�Wq���	�Iq&��!��)�ib�?��#�B{`�w�5��D���Y�%*��DID۶M�R<�3�:�n}y�3]���e�&X�)�|��G��{q&=(�����!Ǝ�Xcb
�]����E��&��{�H�_���?�#0ͤ���u(sd�K1�|r�@q>�
�����~Z�r�Z�T��E�o�\~($[N@9���l=�Q���+��!���)�lD|�a|	��tx��Ì����s�mj�G�C\�����$B�6��k1����!����\���>���IU�CD�����5�?0���}wIj�ge�p��A����ǖq�ޫ�5
���D�����`�?�e9�d�@N+���=1�FF���9h�I�wj2��ܬ꺫6ˡg�/jҟc&!��������������ۼ�r[|��Xkx)����Q��꣞d��Ϊ����ub K�1tI��'��.�W1rtg�O3�8����	���Ck���5�0&����D*]��u5z�`�O?�ľ�Oe8nK��i߫�g��-��$|��؀-���l����@��������0�R�nE���t�m���ӼPs�c�^�h]徰?�5�����x^���=���<t�dS.�f���C�� @+��كq`!J'�fr<\��)��w�V�{����*�|��q���f�di�O=���1�	�~Ƽe~5���ۥ$h����l�O��Z��e���y����ZE�� ��I�:�s"Ob�W8� ��®b�/Bv��E�Ŷ����I]4PhL"ݢ�Ic�,-�g�B{��!o�������X�kU�A}�D���?֔r�Z�i�l�۪�]`�(Q�=�i���/`�i�����r��D�Ah��߉y�`�mm9���^�A9���S^	K������^��r�?R��b�߉����<����H#=;��6��Nwui��B�
��rhLÈ���ӸR���x�rv��_�!bؕ��X:2 h�x�2"�`'�[x�
g��n�n����/|�}�	G<;�;gjB�i[��f�Od)-��{Y}K��|�9	-�13�-���>����oL�_��U�7+�"k�m+�27i���M_kf&��gC��7�Ec�	BDyWKK���<�'��&J�[�Gy�S�zsދQ��<���aZ���½d.�{O�H��=,sm��8��<�"����b"㸚��:���4$V[GS ;���A��1ō�
�/�Bw�11��\���)�+})���2�ɖ4�)4�>$Sc�?Eߎ�X�  lW��L�����|����Ip�m���Kh-�`i��+�(�#%C����1�V&�y*l�.AZl����	�M���}���Z�֖��7������(�H�Y��A���m��/�4�"��&��C��A����8�A{HtF�ɣ	̲�@�*����l�p4��nK#5HC�5R�jq|�n���\ހZ����!ծ�!]P����?C������E&�P�M�h��q	� �I�M��]�͝��C�����Y�����}���_����%�ǽ�TPya�S��L��m��t����*�z��9�b�����LN�t�5L��)py�y�TG⌠{B����
�+w��C�X��U> o=x�t�z���A}��#��ɜ�S�*U3����sj�K�a�����W�4���N��Q�g�)E<���cY
��YW� �i�w��?#����U�o@�'�b�S�iW#r *o��Iy[oFI�D�^N���b�L˦�:�͚P��[W�̭�"�Ag�j�>�uW�ޔ'��WD"g�;�,Ó��Y	-7�	}�n��GS�_h��VP(r�}�z���WdZܼ�X�%���B �Zh��w�D�2��!�O�oͧx��z#�ܺw1A`<�.��ڞv�v][z)�ѨaI��΃���
��N��:m��-Pu��;XFu��!�"���BXK�NC,�+��5s��§�V��L����+��+)�n�3��ҷ�"���a,{Ә��g��L��Y|��v?�<Z��)��=�o�������Ha�} j��Gx��]����\S��W%����(k���iM���	��&����p^�S��b����ʅ�M��ٚ6+iI��⇽������ب�j��A�|�Ț�'��0�8d��Ee�������5w�65��2������	��:2�L<8��>}A��v����=���e���H�k^-�+(7�C�U]�lYO���w�#����l�`<^�`��Er<A�f ɿ�ۣ�T�{^����Ȳ��6]`k��p�Q�{��ުOUq��TxY��D�5��r����q	>�*�B�W H�&�yL�Oc��],Dm���M�<���i{c���p��V�K	A�)�a�3O��7(��J�/p"���6�U/���Q�����"#��[]8fl�^uS��K�89�E=�H�48�8V�D5�o��c?��/�!cĸ:&A�q�{]���)��uS�e��Bb�t�c z$N�:��y-�I'�3�l��s���τ.�|�C��M>��K���r��[���F���u]n�S]�^����׋�n�KX�
_'�$@Y��[�)]GG�D�LB���&��z�K�γ	�j�P}�X���b*��42d�*��I ��F&����I]�v��a���gU��q�^��t�6�����|
�Qf�0`�&��Hi�p�����CvR2� ��M\D5U�m"��"5�`�'�������>g�R;�+iN6�l���G��o{mr�B��{�2,^���F��B��7z�W�*(���eb����㴪M#��f��i���O�(v�ɚ��C1�a�����glS� ���3�K�E6����%��R�]5��@8�'L����� k-�ڴZ�V�%��ط�w�'�9�)Bs���>�̨�	�^b�ƴk0��ǥ�ٗ{�׬fbat�E�#J7G��_�xyq��չ��f�u q���q��	7���t�ԠE�s�"@W�P�\G����W!�����@BH����tz!`�kQ8�Q�1����׶Ȉ�gT>�0�a,��Q0���s4g4�1�7��R�!UdV�;)&��'!/�u�q�D�V����9������y{-yq�XU^'��tvF��B�*K��IB[[��m�O%gV̭��#�(����I�P�����-�0	�� o�x�߫�Z��xX���(��.��X,�R�N�����s�-yaݪU��Yw���+���M�퍃�����(F�0Ex�� ��^�0:�~q��Z�ʐz�yPA�Է�Q��M�9���c;�P�א){u�ƭ$���/��I���l��+�g�m�~��צ�.�c�
[5+�pӡ�Ⱦ��]O���C��ʱ�;\ڜ� �4 ;8l�iNz�f�N���p��y��'���C���`����l�؄�7v�UY�W� �,9�單�tt{S�2�$����ϡql�M�7wpFx{�2�:���^���9h�vc^D�`G�#s�&~�n��������ޢ4�dL=���Hܴ��O�?~�Khv%>��2채�9	����Ƌ�R2��0l���YH��)HH�HD|��h3nW_�[����O��:�m��-V~�2B�2��ֶ4>p�1��ku�G$jJt<Hbny�����fm��ǟ�j;9F�@]9�W�'fĽѫnjYY񃊅�߱�����/���F)�#�ȋ�_���]���{��۷�j*�⧂l2�8����������iO���5��[x�Z��B����3�F1U�T�(`�Qʧ'�Nf�l�݇u����-R{)�½~2O�3���5Bli�nb�#0%7"��)��2C���&����`sġ�}���2���������t��OV4��5�$ne�9}��'O��k`�"��;bئ ]�kڒ�Y��3�N�Tloٌ_8b���b�V��
�1e�7�ޢp�^N����ط�����)[l�Ʀ��E��t�Ǥ�/����ɝ�7@j �:-�{}v�s#|p��m���ĺ��Oe{��S�8��|Z�Uf>����
�X@Pd�|������䂭3�=mb��x��H�r֗�s��g� �.]��ʉ�ڕ����߲p�b�����q@@��5H�J���ap�,�y�����3�!g�.wtG��� +|��Lltن�֟�Xga .%����T7��Ts�8�oG'�t�ίөfOlovY��x�?�J�Jj��}��7_��XLD\��E�B�VI�D�|Ǉa�����*Iȿ �F��U���k�`�`��.���ܽb��ؿ�4��I)����ʋO|����O�9�v���Y����-�̻۩�O�����T�_*�"����1_x��o��VR�D҈��x<���n�
q�d�-,׵��v �mct�2�=#��,�bkbi�-�<�_%�%*���A#�@���&߬P8����X�AT4��xg	���`���\p{� �"w���:��K\���kH���QL�7�����̑����\�#�)��?h~d�h���˞N?L^Fw"�f��,����#�D���1%Z[�ib�pKzkg� ��:k���u�����F�P*0i�k�m��-���=��<ibTb&{~�t7��ai ܹ��0
Rٮ?Ti=��aħ����.m�N!k������vo��+)Zh31�fZT�������R��l�e��<��r��8�k�O	:���r��t�S�m�eeanS5[�B�Bַ\���Ը^���٢��|��5�#o�ޡ��
�W�U��>)�����_F)�}4�M-z�&���0��,�2R�U�2���Y�1�;�KQU#�x�`���d���sbI
S��+���9 �#�.is�b���7\5�Ǵ�<_�E���p�q�@��E�4�Ҧh?�2WZ3�|��^F��v��OJ������
wv�yoNb�n���,<��s�h\0)�-�i�&�]�9����ኊ�~�\^�rӺ�ہ��)D�	���c5�u#�&��W9h��1�{ҴZp�U���ξ*~ۍ�m}�7Z�$�.�-�8��Ŀ���qp�L͹�L��j�_ۊӺ���T�
��W��[�m��:a��y*ǵ�,%���48�����|:Km�e�:�/�A͋��
��D�T�������5Ec��˜�d�T�h���t>f�o�&w�t����KEK���Vp��������[���O^1�9S����Τ@��d;7�.Q���x�@�|D��;�?��5zV��$_xŢ�0ɽ3��Y�xm�5y7>�0N:�U�(�)�0���6�6k�:��F��\=��б�*���� �b�r{��Q � $�09ކ5�]�fR�O>�Ib���_^0�V��T�ދ,��������}nS�)̀ɟ߼.+7���k�;��Y��<tڢ�6<�e*'�\ڕ��>AX�����	SA��ɟ��2�@Ӿ�{WG5�%�IO�_O��=�C��\��/�諏��B�H�|�"WA�G�az�eP��ឞ`�E��\c�����9+�TJ�^�:6/=��!T2{�T>T�j�� ��nj}�Ć`�s#�R)������2���	�=�D�S}{z}��	S����a����J�}�Ա�|�}R^C�`5�[.;�����1�P�m��\007L
�ϻO��w���̟1�md�T>���4�kw�����h���k("Tb��kG[��C�؆�>*�E���s��k)FQ�%i?)��H]����dv��&	�i����J#dw4i�I$ t�tRE��@��YC�S��k�>6�k[>Z5p�p��.� l[9=v/��J�.v���2��9����������H$��SK9<fnR~�c�^B|1�%�r�Ε,�2)��w z2���Ȑ>/O�`��wL�i���[:�L��b7�����
G�]��@�؟����$�Wi[Ʃ4f�jVg���!C<�Zk�`��K!HŏP��.���Ɠb�P]W�z���R*��t`��
?sEh���fVag��������Lv��4����;��M�w6�I�&ە��#W��+��y7�dEJ"8|�:�;��:�z�$� X���i���D�j�`����@�����;]3pxSL�E2(�C��BU��O��KD�Ľk��w峝a�5� ��pĩ�&�a�r�n����l�3(�Bi������Bpc�T�~���^۷]҆��Cm ���*���z�.��C��5�p҆|R���V�;[J�f_R�m�,"��z���3�Qy՛x��ǡ���P��7��L!��T�8��W��&��vw��F%$��sJ�� �`��3ԛ�9��5U�|�C�s��o7w	��Դ��AAP�� ő�w�WyT$�����9�v�����rc�����Q�M��d��Ƕ�����d�pŏ٩�L�y� f�6y�2���bQ�nD7|�G�@�N{�xs�)BV����+!�J͖^B\S�k�,�����twY�Z
Qe��j<�gU^��O7����We�#y)�}������r�h��Z;�
����<��U�����C�J����?_rs &��G�z��|����hf蹷j�se]�=�Q�5eU�+_��L=َ��xZ���P+#�H&7�xd�����o
���+�
����$���.1a�	�,���}OΔ�0Sϸ̭(b���g�Rc@�OJ�_w���և��Q3d�6���~��N��c��(����Uafb�fW��,�CD[�i�l,p_�p��������9��6ꪢ�#�r�6��7��7T8�{�/{�;�ݗ$e�&tEG!�b���iE�±��"�]a����Zِ��G�.d��Zn�1���ᚮR����<U�b�&TǤQ�Ϡ��ʮ����1��A
�)+*�sa"Q��ʽ�M�rJ	,I�d�����p$9fi�bp�}��v/��9�6d<��T�79���yxh�AxwطT�x �߰�{�� �Q�rpV�>W2lc��^�&o�y�[L-o%��3��V�bb	�å��-�5��1��ٓ���1e�F���e��{��Bf-Cyͪ�g�:�6���7���S�V�1s��ݬ��NB���v���F�Z��:���΋H�^�7H4U�˝�@o)K��7U߂m��e���<Z��j*�̞HJ.����#�'��@�^��^+Di�Ou�[8�CFf_x�}m@��N���t�O�v�̿��g+���.ۄ7�]<��ž�^Pc�b�gJ\�w: ���D�]�p�������=TOiG���S�ݓ��Hʓw�M���T��L{�W���Ͼ��} VA$��E�/�����_����\̍�]˫��}a�F��Ҍ���1{��D!�)�L��v�����i��xǘ��U��W~�@�d��ҽ�)aO���"Ɇ�l�0	�ꈨ�2=�h�����Y�^������9zI�a���X)�'��3oG����@N�$��m��Vk�J�ўvH��%��^Y{�����.= �mi����͗�(C�����[U6'IfL֗k /�uР	" ���ӳ�z7��V�H`���;�2��J���	�\�jO1��BQ�w��ҁ�T�ٸz�qn�s�[k�E3��� 1�G�p�?ν�~w�����uu�P�@�Q{~�Q~�@�=�݃�?Ci �u2���}����]j��	WEv\�ٝ��t�I�g�����G4�m�<�Y�x�jZ�ksB�á��Z\�7����NdZ��. UN�n<V�XT��--�h(��\��IW��ֺ2z��� U�uɦQC�0
��}���k#��N-��tDKg��qwH!�dK�M_�=[���K�}z�r���e����䧸k�&O���9�3��f�)�}�;��2��bJ@��y��$��Q���IN8n��i���5 ���vH�)ȵö�εA��枳�4�U{/���3��9�E=%��h��zu�*3%%G������.���?*�4h:3ʹ�K'�>ah�e�Q�7@�pbϪ��9q&ι�1���^��[�BV3;ç�����]����إS�f�a򔤁�҃�� ����ݫT'h{xm��y;����ӠhL��Drqg��462��*u�`O�dNSʐ�!���+"<��G�6o��>|�vA$�&���{�]a�)�
�'�g�{̸�xaHn���$:�5d�W���kVW5�wl��N��N?�^��lj�AW�C�Q�c�7��}�3�����Ҵ��8E��BI~%��w_lڦAR$�����$��­eB��>s*5n$G��{M�k������A�e���Y���L�9��Q���5�$���.��d �\�ll�����Q�"�xn���}�bB��Ѓ��fV7q9�Ã@ <|Q%���H��'ǩ�/����.d#2PU�x��ۖ��viGʺ�$O��X�:��/�gA��.r�����`\�����]�-�S{W�5e�fz�$��O�kӉ+!�c�T�}�'�G��B--��������٭�V6O=i�r��D��{ �m���r4���&��j/E)eNZ�$v�i��5 ������E˅�\$c#{��|d�0�Չ@�D�Zn98)h�aD%0�����#)9瓕���#����7D�Op��=��;B3��5���Dt |K�e�P��)��*Z�v�;\
M
����;3;t� p O����7�&UJ����>�yK�c"j���ёK N��>+���S{J�3?j.gu&(Q�w�Ю������ �o�N��l�ǄK���
�zA<��?M.�{Ūj�}��f�i�X�y,MW*oDly�g�PDt��I0D����xh�%��T5�,��Mb1C5p}�����|{s\\9�]���kzA�>0媋������I��lÜpAꍟ�F������|^��!1h~o��Y���7$��%o�ś����
D�d�����I�<Q�9Ua����n`�[c#R4h4����6���b����ѳ����׫ω i�5X���0��_�ѧ�%X�`?uJ�TU�χg�n�*�����h[��
;�����`�Lbu�q�4Av�����:�4��P}<����x�==�����y������X���o��`9_ZM�I;��m���C"�7d�j���?�E�s�(h����8<]t�2<~Įpv��6*e�:ם�7� k�5Mz�֜u���0hE>�`�� S�t��m#t��j�����v����:������r��0EBm�,�J����iA6Zݸ3�g���:/��a#��Ŭ`�߱>&��%��g�rZ�*��H��uU�`����	�;�2��e�P�XÁ2����NQY���u��}�Ir���ʏUY��ى8.Ӽ.�s�G�y��؜��mr�7�!i��� ��k�y@"�Xv iv������x�_tA6WyҝmM�o��->�ed��Z#�[`�A�c��y��Dy�ҫ̂�v����@�#�[[��h ��7�&�)��a�j�Gc��R��i,A:>N�<i��fD��j��5U1��3W�hV�Vʲ�{��������$����VZ����Ϸ�1b��MM��N��#ڤ:ka���Z��3��c����z�^�~��GS���dl (�T�Sl�_�&��5�7$E�??J���j���W�Ñ0N��I��r�rp1$�0�9-��R�	b�7��zQ��H �kn��ĀdI��Ѯu˜��g�8��I�,PJ����	l@��}0S�M����|x��s��<P�l&�Xrs5T~35�����6��Ea��,8�zv"\��8��J����H�ԟ���������knsbb����~ĩh��)k��r�$J�_����bU������p,O�"_�g͟�$`�G�Nd�'@g��;��z�v�����	i���Ӌ��G�(�ߠw�%�'Ж� T�Xk7]!E�B}����h�>�!y���<P21�9�6z#��#̆@�w_�Mq�7~_��t��o��}
W��y����YǴ]Z���l)X�8��G���jF��qS�]#�V�ă 5�'%� W��v��[ǁ����W�	���ƥ����h�gO�C<�����b�)�-�N �zd0E\�R��O�:ǆm:��M�#��?�s�|��SvYF�K�3�k�bd_���:v;�f��:���J��M�^)T$���Q�����-���y}k\�&f���G���,�µS�x�����1r�����<�p t��`'���u �����]|_���H �;�\�8&��Ŋ�5y�,7�Q�r%��`�������S�[ =fUҚ`/�ξ�۵qܒT����|��?��	��Ý��y�+cL�z���� u�TV���e���K�F��z���XU
Nt�=�$2rA�5�9�7�(܎�i��(��q=��.�$�h���m���`��:�w��ܪ������9ZX����/'񩫖�ş�<ءg�Qj����Қ+}�L\�6<�^?1���r+��Jk�5��V��p�Y
�4�u��^��ӏ�|a�+6�*����[M�;��˅>GZL~h]m�l�s�J��ӓN�h'��k����
����˕�a_^��=�z�q=����� 0�.������2�"O�uX�Q��9X`��r�ΙW>�d%YS�Z�H�\�b6�=��1/��ڿQ�Fm{��rr����d���Ϲ|=�*-/c������tߋC�/~^��o�ߥΦ�I�Xٞ�����;�.�{-GP��C�ӕ�%֭3�ߛF�`
N5��l�.]3���{6i^EW��H�S_���]��*��2�I���"�=%�"-fT�^ (ϫ�ޕ�*m��h��/���#�e������o�Nl$С%ǟ�W�~���|�MChߞ��pKAX;O�~w%���F�� �"D�|���[�~��?��ÕoMGQ�9��� �(�9���Mg�3�M�J�;�2��'w�9 �(���m�آ�t��U�i^�9�����Ro��)�p�������9o2�Cb��1�\F?;!
-��k�Is)�OɴqT�
Z���3�ۋU����� U��>�
�z��ڔ�g�i<Kp�����=����	�� ��K0ebUsj�y���!���JxT�_���&.m-�����X>��~al�p���xW'6xL#�AGS+N�"�� ��afb��,�� ~:�V:��n��e��|S[1���ʋ���㧓��5�W/��k(� IS�Z5��-[8�f�$%zw�9�G?�p+|Вz�P���o���qx�r����Xe�����41d��Mj�QO�㲪���^h�������$�ԊJ3q�2ъ�c��j�Id��xwOk����W.feN���?�ۿ�i�؏Q�N����\n���XSM�`E��lM��-�6X��<������c�H�H
��a���&
&fG��
S2;��7�_���d4}IW�_��ƹe.�,!��������`�^!0�O��ſT���G�� n*58��St�����wS��K�D�/~��&���,�a7�=`��/�l�^�7v�<�v��C���;��|�ў嚃e��+�p�QD��yQ_�Pf�"���fދ�99f��Н�6�9ap�r������-��Lid��%��i�*�N�H�A�sqq�W��}�U�}޶��'��p�[����;Q�Vٳ�	�l�H����YQ�-3��C��p��k�W�#LjЯ����b�<��aVЛ�Y�IJk���U�e�������x��ڻ2zR��2�Ӧ��y:�e�<x5J���Ju����.b��J�����zseuq���#��%w��Z��R�J����/"X�ٮ�޺���s�_J�vl̚�c�c<���ر΋�܅�mO{z��N�n��9)2ͮ�:�)�l���Ǌ%��j���؂�BPƒ�6y��g�d�a<$"p��`���$j�q��-�r��H<m�̭�\S�'.P���	J$�K�󉒻�b�Q�)C�4���q����ޯ)&���q�-�|�3�lL���W�<'���Z�&s_б`��	6�=*��V�(w���,�M��F��C �'����:��:�c��2Oq{�g��N��@&�S��\N�����J>T�QFvt�R�7����!#��B��ϋX�|0�m��Koi�Qu����?g�L��r������ɈI�t��\u'��6���
�$�0�Qe��r��qSԍ8sJ�b��2ln����Q_�;�,�#%�[�CX�񃛔��t�� >�*m-~4P�hFۓV.2e��~o_��Y�Ke_�§��׎�>��XZ��s5��L���,��.�P���a**�i�w/���ޗ�q�m��]��@��$ukҁh�����Dcٹ.f1nzdQp�ğ&� WFjI���W�l��+����g/���=��G6�9�^�J��(�9Wͩ�mlW����%ӣ�q��6��:��H�q��+�bJ��j�W�Q���p?��hqgW�����u��.�{��탑V?�˷8��ƻ�����rf^͛������m���X��8�����\bI�/���4sz�������x]q,k���=֫D���g�E?��Bj[���p˝�Y
������i���z��qB�n�b��I ����oU�9����l�hR���L�Xll'F��߅���k�r�L ǤH�V��vQ�g�7$ƹeq4c��x�����[Dj�Vqh��#��&Cm��X(��à؅�GͼE��"�\���U�.=q��Q(�z1}���j�<^�H���{�#l�,�w�4�fz�C���3�%����bW̍���T&�����H�3|�r�M����i=�J�Oa\���PyBv�ϭsa �P"!�˚ZA�����}c����L���A ���=�������^Oyd(n�J��p-��ha���h
����j�6	d�5�0�;#a��ε+� 
 ��W��pu��?�\L��
��rJu5+�7(*) FP�؟�h��W�k��룏6���ן���-�f�9�%"?�Zs��:�1/���N]�C>w�-���	�h=U/zJ;� �Z9+�l\��I�0�3�zp�$���ު"�ݮ������w���SyO��g�b���~�]�^]�+.s_⏼p}�RHv�N��(�Fr>넵��(�����A/�"& �p��kl�0/��c�T�E�V��>_}�SYH�tJ�w�4��R��.
����P�j���p�x.j�_C^�Mm�AGz�$���=��9�n��YMW��aP�5?��Q����Q6j��9(����I�{R�O�`�����>�Od���Kg�92մț�9��Ӷ�0�W��t2�]̚L��9V�Z�y��@Taz0i�GG ��ɩ8.P�oKp&�(=��`8-��0��q�,�1+�P9������p���[Ӄ3g$���Z��q��ʁi#��N�j�R~�ͥ��$�����[���E(�q6�{S�|�?���Ҭ�:'��=ȕ5��-hQ2nⅸ#�v=���5�Y��{����<}�Ɛ%� ���#d���C)���}��{��xi�m--��1�X�T�.���+ܿO���C�@�Ӳ�,]���;���Wð8S_��j=3`�Ll��ƜD�Ǆ�E�-�&˃�e�֑O��k�W.�,��	OL�)UZ��u��]�L�|���wL})���d+��S����%�J��&��c1��	��U��H��lskt�j��X6����
g0�Ä:�)g�~�:�.;�ט���e6}B�z[�?I$/������ R.��aדq�]C�+� )�ͣ��&{�Sws��%@%3�������Q���% � ׿�z�w����;?��|��P�`&�
�Z���B��"��?줎��cn歠���"o�g��	u�P�_R6�5xŨ��v�a=l+J��~�}?(�3(�ZD���K��K�Y�j[�Y�����~V�G%�7<cVj!_���5I�@�3gS3���;o-�Y��S��w�Н�l�v���S�y�#�����).J��)�p��9��.{0 #>t�q)T
��7[cr,��W�[s�D��% ��r+�����x��%Qy5/R:�^��1ғ���".��l�3�zbO��}1�R�Wn¢$7�Q'Z�Y-&P�յB�O�.��*ߵ�l�`���%�l[^�g�B�rõi����Q�;�{�V��챝��l�. �c���-�X�מ;��.5  I��Ir8�4N|;=���N��ŏ�H�Ug�q�(�o �iΚ��j�M*�#���PaC�@e2}t�)ŶH��t���d�j]^�d��u8.�-�,q���F��x�i_�L�p�h�L�q *�{.v5����s�<^7�)�sk1��(�]����f� Ċ{���kP��OZ0�Tt}�9����/q�`���R���\NȠ����K�=�Uoqu��y7��55��q�:B�m��V�|�@��� ��z�(')<+Fk���b��Xĕ���ɇ��I�4���f��E��8�fT�����	��x5«K����Qe�Z�W���6�U��n�3�]<�}a<C���~���(��"�-N�[]�e�"i�D�����i�L��}5A[3T#���3j�=�PJ�3aa�Yym�Ry�ԃG�!�	KKM;'���nͣ�x���Ī,I��>c%��v|���䣣	���OJ8Yז}[h�n�tX�V�<�A�牔�X]�.��F��@c+`���HO�y�&U.lX���|a�A�a�Aޒ���%1��v�@���V�_���i�z�^z�eI�6s�VxW�-��2�^�c�O�$0�^(V���?y�lm�u��0Y	6�K����rI]V;z��0�a�e�Ѷ�Ը�	Ln�>~�ψIM�_2���5M�ДǇL�B�ȺZ�O��V!$:��&hg�����cG)��aL%�*g�mC�dcY%'���yl\�h���T�� LāJ=VȋD�|���i��7�.�I�G�&G�D�IK R�r%Y�9���Y�v>/HW��*o*�9g[t '@��$q�E	<��J�R�I�ٵg��*d�3,H	-C1=��$f~���0[��UB�Hd	1�� ��(�9��>X��y��|�NE-����n2Չ�z�tgb�,�ڳ�!Hɨ���̀l�����[�*�#��|EO�D�A�rLM�?φ5G�1���W�e����j�TJ�!�C�e�'���"x����K[vQ�5TY,�M�q>��m��?�#>�]�wvX��<+�v���4p��� ڞ��D�F��\�K�|�����1���e������FM8nV���Gszf�W�!6(<P����}F��v�T唠��_�N'�i�^��Q��_�%��[(,4�M�MW���>�+�н�Nݪ��n�U�%i�����L�-�����ڶ��{_�� g�֗/����YƘg&%S��I�UA�@����ۿE�"e.��C4F�{���>�����A���H��G$r~y�x�-h�/���9���è�1ܽ
�Yu�c��S{X����*=��4:B�F4�����s�Rn���d���u������1l�0(ty�-�Ms�şfE�W_(�eXc���B���.�dfO"�R�g�Y��`�g6������ę�2ُP��̾'U��V�� 0�Z~[%��C]n2� ����(��C5�[D<��ퟨx���#��	f<^n��t�n�
�s��h� �IL�Sn�}�s��D���������W@XFC�&~(��5/��P�s��y	WW�8�f ��4}CM������@�k^�EvH�"Vc�\��$
�J��ĩy���
+C`:���&��M�=�y���J����q�����n��BU�P��( L2�y����&44uۣ��+l{ꮟCݯ���Y��͵I�?��o�p_{E��u��w,�&l�4M�B,��mD�����C�Fw�H��G�nr@��{Q��\���`װ*�f�T��e�lx0�Yyi�:ˤ.���Z�\�Q���Z�U��^�˯GS4�5����oK�)i�u����C���)�d���D�/��R�*�&/��_��7&j�� #e�������R[ɰz�A�n�	1��H�>B�LJN�����T��c�N�C}�F�<mtC}H��ר�G�����y9j�|٦C��3����������r_�Z�%"� ���(��l���4�>��eHm�k��~K�8����m<̇���*��*p+�&��G��Hp��Kan8�=�g��-��/�|�����GWː��b�������`����we%�0�|��o!���/�YD����9��k�Nb<��& ��}��}y�̊���}f������)��#To�"Ĭ�G^�n�
sۥh��2/��{���Z��i?��҂�O�8�5��7]ML0�'cƵ�����_�y��sz�R(I>ʕ��!�ћ�&�J���5���`���OѾ��a��*��m03ӯ��n��%�<x�'�̛��Nk� �.*X�N]$�W|����`�ܕE7ˊ�:t\�nt��{L�Z��5�L��+�"�7�%/�jg�l�'ϥ������:E�K�n�>�DCӡ5Q�s�
��aNAX�
H2�ɳ���ٱq��2\��E���PA&o�[f>�M'�#���wo�?�y���j��7��{mf�U����`�ǘ9�;%r�p�����˯��J�C�?��>&;H�P����ן��{7`����U�5��f1�:�	!ڰ`�i����<�c�F���B�M�b��A_�4ǬV�P�U}�$�kF�K[5a&�*ݜ؀2��Rx˺N�����DE�x��X�d~/*%�#���2b��Y�6��{��G/%���Rx��_q���,|���Mq����~ƕD�;��H#�'K����+t��Q�aXb��9��+����"Cx0Ak��7������j�o��jj�a3�6o���a.J����m ;3=�k�t)�	:�9�{:T��8{�ڭCK ��t_�S���v0�����m�'����I2�6LN��~�#\��o��4ZVH�}�M�pR2=�s(4�0�ry���f��Z�}:L����������j����3rY���qfݺP\���:I��tɖ��}�R�=!컔r/�F� ��q4�Lŏ�Vf;�*i��̉8؟-�������	�eJ�jpR��G�o��h家-����%T��	�$���8*t�~���FPG�@U�ፓJ��o�%zb�<�C��ಕ~y�+
ћð�`Z'����R�a�,��%מ����^t��*���?v'���o�
SԤ���ګQSJf�q��
tq�nb�:�&�D�7̈́�Y�Tr���"�5��'25�$�O����&�b*=��@Y?_�-�&��vj��.3��4n��e�[L��ux��"@��umQ�ɰ>�nU!�����jD��e˫=2��4E�J�&��v�z�*]��N������v��7��u����Ζ6B�ͪH[T,�f0z4�GX�M'��*?��y����/m���h�`��_��;���y�Ή࿼n��:*�)�d+Z�L�Qz�fll{������@յ��F�q���	*�9_�Z|�cx��k6�8K(8yu�f��Ue�!B�NJ4~��+�ڹ�n<����'D��?D���Cw�y����M�4x��4�W�PÔ�F����P�)?��GmL�(	j�,��l=��Ċ��k�Ƌ���_�y��+��>i-�B����Q��*�G���
��F�ӋE���q��k����N����P�J`�i��U���+�_"�&�4_�?r�Q6bk�~�:����O�S.�\.�+�x�@;�/��*�<X�ޯ��K̇���U	X�*���������8;��B�(Y�M*�S�o��>�5�#��� �t/x� �DE­3)Q��0�7�i�f;��q؇_��!���?x���;�В�!_5��P2|1�����TH8�ē0-k;��S.�w�=���g��S�X��p.]�e&e�RS��G�E�])mQ����S3]�V� �{�(i�>k����.���:ˬB�@o�<�� ��-G�`�?����}��2�CF<�9K�C�EF�*
��M��Z�u
`����A"J.1���Ut�~9,�gz�bn���9dv�lR�旙�l�/Ҽ��X�Т��AXi��u���w%�;���'��j��A����
�^g�w�L���>:�W͘�nR�����2U&�{��Sohkƹ��GN�����/�0�S�ٴ��bs͎\鲤��Ɉ��W�%� ~et��T�^�ܻ�M,A��W�I0_I�PأFท"�uǀ�+`�{A�rL,-�OG
n���9��ʻF��	��O���j�n	�1�i��d�r�!�K�@"�����i�rs��x����P@'��'�Ge�$G�\h�U���M���y��y6I!�;U��̟8.��5�jA��A||����vaS�=)~�]ʣ��=Ud�}8^�x���t��"�6YM�۷8Βh�����m&�D*},��R��?�EJ�1S���	;%��C�l�����e/��G�>1O��iU�w�b�Q������-�͒��%�)E�%���^�旌S?�;1�9k��L�E��!}QQP!����?��M�\?�73�;����@�́;v�«
VH6�ڻX2P�\�`ﲹW��t��M��m(����%���5�FM�C�?���~偖�Z��h�;�vt��b_�,�m~������X�鰹uj?�j���?�q���(nU�Α{(F������{���}��Ԙ�_��jkވ���-Im#��I���z�-�T��G\uN�#��cS�>A7�������z�5}s�}40�����2�N,p4wnV��`�a}*h��l�11TN���ܴ
s���oj��\�����ceTd���;���1��o\�O+8�KWn���ʥ�y��~��k;�J�W��f�&\7r�!`q���%$������t��f���������)G'h��zcNL�������)�&.�'�������f���,�G���#e_h:Ί2�Á1R�B��d�]s�J�U�������
%Ōā�`Xl��n�[x�c�a^��Y���<�C[�Oմ�:��!a%�j�!��7�0��T��A��g�'��K+�T3[�}:\pϘ����.�ywF�
��	z.|\�/(	8x��v<5��(�N����R��� ]��7H��ٜ&ٮ	_غ��q�)�i���ڥТ뾐��03��h��0��@^�I�l�f�f��\|�»�fy���JN�m��
�ϲ��� �(~�4�M�=�FO�t��E��e��}��g��Z��b�gve'}8Ae�UO6�Y;,���Q̭������F����O�S�MK�1��ߡ�iɐ9�@��~�v �7A��2�&��}b!��2�肣�S�Co��zHf?����է�zT'�����Ť�b�0�%Tq�M�Ef��$���x��S��v]W�prl�I��O4b8f �R�/p��1�-�h���S�A_����p?�%��o.vO�Q3PFD�ű���+��E�W��(�t!ދy�:���1Z4�rڨY�z����\Kch`�,Y�����N��!׺O��!���JK��J��O�uE ]�#,R�t~��hn=@(�ʻ�}�_����b��p-9sW9�������u�t��x������zY�'����=����h�y)�=� %Q/S �j9�͒I�c��6��/W��/��wi��4�f+�v��V���*Gt| ��X�������Ej�G�Q�����0$i?��	$jx�{/=����]�2�j�F�U��	�~:;`�3�08>N��ǝ_&�U���7y	YT��9�Q�b`%ulG�Z�pGl����*oP�oeL_e�j�dw���U�~��+$r��6%�Yx�B�>Pe�s6|�U���wi`{QW�NHQ����T�!W@u?�;��2]V�`ѵ�_f��8g�w�-2���cܨF䮊M�W֧k{���U�*Ao-Ѱ�N�.&��L�D�z��?��:*R�*S��>b��l�w��qhA�!��n��W?D��t��J&�f�5��,,tA"�v�z'��v|0���
�`b�?`zBm���,�<�vwl�R�¶������"r�g^��^\Ԛ����*�o��[�Ѝ��+�KH�a�2��k����j�;S62���C�6<��FL6P��#wzŷ/�9�bP�,r3�u��%ܚ��yyP���Ε�G8�#�{�y�%`p�9Ov�b)֕�Y�x��*ՙ�I���$i�⤘\�Pc1X%��H�7�la*耱�Wq�eY��{O���5����[o���e�/��^��BMU־}��e���`N7�ajA�(ׄ:0f Ho��UFR��qq�<�y[�=��^\��a��!9�F }��T3{�Z�z�HDI6�,�}~�}�qD�zj�Ǿد�fP�Iz��#���beM�jI�������f,�Z������v�ڒd��S ���+k�	����G/4Mj�5+�s��Om2��B.dU�{��كk����D!�s�"_<ͯ���TM�6˺	�i>Hz,��W9M�ɘ1,�B��]��쇊��/���UA���{��x�,��c*���0b�t\�T�#�f���lK��-�i��V±�ɇ+ﺹ�*P'��f�%��GD��r�}Ӡ��k��.��4�L��5��ip�z�G�e��fl�T ��N��Yj��de�KO�E�F{=1�J7��I>��^h��b�g۴qN�=zѷH�)�Y��W��-g)�f�a�pG�������w����r~v�B'�;H�j�$D:F]?,����T�z
:>1/E��Q?�,���7��F=i�@�/k���O�@�T-��׏WN�������Lia�b_��8�+& �D��l=a{�<TY�-��ߤ�L���^��bOu�
���Žo���ރ��և���!
��(5���c�g%�e-��$D�����-ͧ�ȣJ���җ��@z��<_o{z�ړ�p��]o��<,o�\(�� ��&�b�@A ��\��Ŋ���T�K����|X�YB���iY$.����u7:��wj�}[��	<e���9*#K�I���q,��K�v/���� ��FH4�����ɂ�k�%�{n��N�Y�f�
�;�e�68���8�`��[c|��GE��ȒJW ^��Q�פ\ꇵ���@�L�qR.�b:��t�^�������u�0 \[x���z�a�����m�	�IQ���E�c$���{�0خ�/]�=z(t�B3�|���R%�@��pY�ę���E�A��@�5����$�G�ǙK��aR:O�����Ӥ���TɌ�U���[��&��V�1���U�Zq�:$Ise��X���Y��m�-�G5mD��ih���0ܹPf��G�l�G"�]A��ݼ���M ڭ9w�u=`H_����P
O���̬��x,}�S�*2D��37[���6����0����&���t	��5����0����'�������� �����T�t�p�1ܬ��i2	�u3�~����ÕV$�E|y�h�^��68P����R�oG�m�zW��#GC�T=t���J%��pg`���F�݋��3��?d���҈$�����l�PI�D�O=�uOi"%��@)�xŔF-�em�xS|�]��]�)�"Y�8g=��q��>����6����1K�	I$PVM �^u�Nf��;Pe��,�W�֓��ہ+("��צ	Xg� )�.�����\�����X�m�gO�n�`)�܆C#�	��S��$1uEމ	m	��+���B��&��W�^z��3�	�������>듾��׍gM�\3�F�\��jW�����r�
�a�U��c���͠�t��_� `aU��{Āzr[�P;.�Q�Wy0'2 ��&a�������/���$��!�/d����l�X�.�ݟX��8�ۿ�
���(�bJ"�1�W����s��8�h������ W��s{-1)�(�l��t��:$5q�bv0svd��&b2��.:Â3>P��}
;3ML��Ͷ�����8Z�P�{1�O�	Ҟ
�G��i֦�>��J�"ʌ®�Y��_N��k�����Zs��~�O�A���%�U0��KaP�V�D~'���u�v�|r-�iX�}n�}HRI�N
;�������⌯��66W�0�U�A+�]��a>�E��?�'FDǁ2����3Ӿ.R�� �\"���D�
!��%�\&	�����h�27R4%6��!�]��8�����d�L
��ÉL;�}U�2�Q}�}�7�~+:���9w"�={���^b�_}�Ţ������9Q�G�R�~O�I3��C�`R8����ȳ��ڌ=-p���Ы�5|��j7�4,�.IM|<����}���\,�7?УΘ��h� U-޴3������/���A\"X�
V+X��5���N)������l8����8R�$�_~s�v��$K{�H�Oz^\�g�=6G>t�)U���v����aޢ�B�ՃR1�qlTGAO,^�i�,A��}G�8-���FUS�ؽ���8A�2�,���i$hD<װ�G�PU[��w���C�#E[�y�@�qz�'�J�@���Y�#p|�DS���M�9=�ٻ�VB����-��������:X-��j� W<@n�c�͙. �@D	~L�X��prd�k*�|R��8�?ſ�� U��g���т�oy�eC�4`�~ԺE�i�>�4�G�U܀��o���N�����H8���lZ6X��� ��<��A:7��=��q��I��%�O�x��o F������{r�8]�aT)��D>�ƽ�����X6��k*�jS�\Q�'�8V���΅���4R��b��)V�����__f�̲_��cY7]�_J��\Ok" �*��qϺ�5DvJ��+��+?��w'�5���w8���1�c�!`:�u�qN7G�:�8��w�:=}"�O:�8_�6��Ʀ��W�.������p����"ƚ���|�D.�{�!�.y��aWa��	+`I�A�<;?+h��}x�u"jv�+p0ɕOV�>��́�x�,*��{(��(x���ٸ��5>h���K�1��'*��@�(&=)`(��1ϲ<+
��J�SBp�Fg���Y0�X�
W����;�ezF����N��B_�K$@��>�,%��Dq��^"k����\�E�6��9��<�?�b�P��Um5;�%S����.Gh[��#�mXvy�k�N����w0��]6�K5���߹m��"#�G�� �G�E\8>�Q-���aڮ�������YiÐ\��ؕOgz�*����K�z�ő��IϪ�u�H�l~U�Udg���+}	l����3d�����[/4�����eU�v���z
�����&U|�Q�"��� ��]r�>giI��]��q�������j�SتGt��[��h\ f ��ezS�K���vdQ�������@qOQ�8���*��I���O�!�ƀ��sU}ɦd��j�h$H�v�*��Mָ"􂞽U�ԌY-&$��g�Z���8�)?]@P�j���2`ۖ��c�/�٫���\<ܗ�Y���r)�!)ŉE-�7z�{����8¨�� �@��r����t3��B�!!��?����Is�&�{��>�DS�ߘr�F�"@���Y�L��ǛT�g1eJ�{Z͇}l	�u��}"�7��B ;�iWȀO�x�2���N1Y��d`>xv��`��g�r�M7�og:l�fT���x-�]k'֦[�����HX�{.G��N�D�[��/�	
�3���"lS��a����ulƎ��cd�Rm��Qgq�G�Eo��>�4Q2A�z�<��^��r�t������	.�q���������x�S��L;�gG�]��xAo���l�/����/�0��N}BUv>G��
���P�L��q�r��8�C��O*m:�iK9���ʞ|��>��E��A�L� �@Y��R�U��F}$� ��(RB����\D?=���~���E�p4�ǳЎ�o���A]���@ρ���R��?�g@h�19@Yڈ#S����V(X)ƝPҲ�!	X'őUA�d�k2���AA�E�~�,7�1��	բ 4�#C���9��\�扉#w�j�͗RV�o�����H��Z1F�z� y�q�Ei�+���u6��\-Sʇ���̓)\�\��&���'Yaz������|��Xa�(�>��:o�X�G�Ma��������bڥ+h��v�2���[�G�Pd�5q�F��zu�%�P�\�"[c�x�
�:�'���R��^����Hpj�8���i�}H���)b�r{}�����jb_�mh�4���&�O�=��.���!ɄU�8�+9�=��x�%Ў RS�.khU�j':mK�.N���@T��v�l�N'�d��`���ט�g��>��W���dz5Y�%�ӌy�<�.ي����-�)*�U,�2����S2̨.�ףR�dof�}�8X3X@�F[n�sRN��A��%MݛQ����[��)�P�Ѳʿ2��=��Hgv$a|^N�T��C\��=���,����D� \C�m��e�xE�NEsh��CE����Y�Yo�?`�:��K�]r����V��r�֊��c�{�I}�՜�$w�9$�ᭋ�<ܽ���znVy�Ysw��2����&/�+��� $�v�t�@_��bJmQ���u:]B	Q��:r��~C~�����Oσ���6nm��F���M.HQ�@�ߵ[d�A��O�D0+��|���ӹX���q�w/>_���gٷ ��0��Pͮj���mkT0���d~S�u��q)���{�E����&��$��� OJ[�x���8�ԫ6@R�Ǩ��[�i�M�G_��NR��p���W���Lg�ZsO�dcU�6�*�K7]��3r��I���J��;�Y��yUdk��~�ku9>�FX�*zt�/��]Q'srμM�eB����$2��|���?��\91�l��e=9;^BNI�X�6��������O�i�p�'��oY��� =(5}Y�B�O �B���֓�&��}I�(dB��Z���C�tZ 7q*r�ǁ�n��'|��A��5b������Z�+_�ǬQ�.EeN)�7*���S�<���Ny����<�;`^OF/��ӳ;���a3��v�a��a�����	��-	����v���sfFkd��f:��c�H�!k;R�5�#2�r<�5Hh:V�ZU�ll������`�鑥O��N\�N�[�R +�l�@ ��y��cc�Z=��YD��R�n�ۋ07���n�u�91��ݠ&��-D���S�?��A�p	@�ħM��2�xEfU�R��ϮJ9�32jw���#�LϹr�W�;����e�+<��O�ԭ�.��` �?�ɷ��I/a9�^qX���s�{��f���-tW��R���7���T��N���v�T��D �y4}ʽ)�@��v��h����B�_i�#<߷����	�C?���o�������wB:=T�av�ָN��ө����<Uf�7���x_�]��Tԅ&8
H4Krb'����=���U$D��_:8���D�����x�i�J+�#k���a��b󮒳�̭X�=߶����4�kxb�4 �t{1�۞�L`~�\ii�f��fd��޲?�3��-���],7*�70^����E���t��C g�J�]���	1b<#�[��JK*�x�K8ݥ���1/T��_�3zu-�"��p�L��Vƫk��l��� �(�/맅3{��t�5?-���lU�)�g�24\��M��U*P(AXq�u��>W�����B#l�}�t`�qy�B�b"��ԝ{���D���>�$.d-��<�u�E ���{�Ǘ�ȝs��Đ��Z;���)	�,�\�4���ZsR���b���y�=�ȰK���c���q�FYւWqo�[JB&�
���Y@^��Ǜ���1�˦Z��r�e��FV�v�\��Ўf+� �v�E��4E��(\�sG��}�gU&�ي���z��4�l��|���w���C�K�/d�2���3��	��9e�R������wz�������-u��s�k�on\����!!!v�F�~�x([	��З��E.�*�JM`%�Qs���f� :VhJ>�o9yا���Lĝ����T�~DV9!?�� �G��ۢҿ����p X�<�������;�sC�9��D����7QXD��a��5�����?s���tV"�2�qg�n��R�93�7������]�Ykp>Ui� �\�o�3ȥۧ�ux��uu���M�ׁ���О�����L��_*��@t�!t���!��F7��q��� f��ɴ�z��]���i��έ���ȯ��ay��SCdO�r������p�L,<�IZ<��;�w��x����%��9�A%O��QD�L�
d�l��4�Z}]q�9�����a^r��D��%q���<�:	�1a[�8�[.yn>3ð��I|P�$P���C��k��!-��ѫ�8-D�cI4��7yؽ�"�-��Z����J�vQX�l���w(#�C|�ҕ@m�2L�&.��_L��F�gY!`�-�%;�?�d,	�I��������r���x��C?�i�Lz��.�m���8��s]�Ms�Ex�����f�������<�u��LCC�m���܎���M��^j�j飕>k�!8S-|�|�9m���}ţ���τ�'�F
 HvY)'
6�I�@�[�����U����M��S��8%sN�C5��e��FA�%������QO��a��At�Y}}����s2t������ٿ�z��YK�4/��3X?�����Z�R��'d F�g|�^���2�ڵZ�#3���X��0�8=�=�I5�m���|Gw�$&��檟���꟱�F@���;6�s���g��#|#�{�KG�U%���+ş��	RXvd݌l(	Nv���Ƌ"�!Pe�������J`�v0�{G�ב4_+�L++���s�g?��(L��aӂ�W���Lz����L9i&�H��	�Te�{��f\`��?�I(�{�膞��Gi��А�����vh7�c���æ��X�\��#-E�0O
�7(�& �+��N�2dU�k��$EE��G=�'����C��8�v|ӻ�_	|���
b�KNٽ��o�Ԧ���� ��"����|?'W������'�N�^��T��?d�<ְ�A����� ������ƅ"��@�'�q7����b���NSM�*���w�2[�,�r�E��:�u!#5���̲&ת�?�G�*<���g\���{`W��O�s�M��y�=��9Y1���/�f�� {�])p�4��R���qȫe�����;�0�Us$��t|σ6�@��~�C��$ʟ��+�kR��{�)<��Z���ց��X���ǒ~u��؟C�E7�����$����� ��]��#�= �X������69������̐�����Y�'6N�t N6A�]���U�D[7&�d3�����R�1EK�1]��O��{��������,פ|�9�*Bd�¯��E �'�`�G�#�����ؓ0�!�� �2���ߔN0��^�X��)\fJ�e�4���I+s����e%�#61��Bw�
L"�N�Z����R�~+>�yz�;#,�V�E��і�顾��ͪ��Tb�6?���I�X��:Qპ�存�u�*~�n��� �}�Q'|}W��
����l����%�`>�D���"Y��s�n�Ob����(�:���*�Zp�jT�IL4ba'��;G�F�S�$��(�߭�enmÑ7x���e�A�*6�ܙ��f�_z�lAA����pp�j~³�r9Ll"��ˈ
TՆv�	�ҷՉ6��n��N:앟n���V�o-�ΕA$7�.�<���,�Ilߟ��P�?62,�,2�ME��������P�Z�z<v�
f��RsF}x���m�E����u��΋1^J�T��wP����
�d��)>�w�k%(���9
	�;�[z�'����t�!���4���,�_wݲ�.�'��1�߾�o��5�ڑD% 6���l����n��������f?�����\���a�10���e�q�\SX�u�Y���B�5��������Y��z)y�C��#�H��:ӧo���!	�bj\h��[^^��F;�O�� �-X���(J�?s�~��(-ֈ�Tҕ�}0C��Q2*"C"W4�
���[��$I;wpA�<(��o�r����0ы�1�& ��C5~��%Y��VD�H���QI�Ѻ��<��\8x�%9mC�����!$��7��Zl���5!��{�q�'�>�Rݸ�:C��`"v�e�Eh��B��_�4A!Y�˷�!��x<��1�alWY�F�ɿ��r����2Nxp�ܵ�{i�=R5��;�]9yH�+[�=�;�ވ�@�CY�B�K=�6.���[�qY|?O&���Õ�o��#\�4�_��_"Ư��� �a�'�s�خ�85�H�&툞a���2���B��퐈�_8���@�`�6���Ű1��,��a�1t}�wA�� V�]� c�ҹm��Ǔɾ�&fa!5o�A֕Or��+t�uޞbK�$g�R��-Y�߈
�1Fi'=_�ZVB<+T{C.�F+X���/�w���Nc��]E��E�3��g�8M�Mf=� ���;B��)ʟ��Rd�`y
J�D�(��y���{�S�@��9J�$�wh��O���q��Q-�w��g��
*zt�]{���d5Z�|'lM0�^�l�}Ry�����I���E��;� �.z��n&�����c�gH�u]�7u�ȑ#4r8����N(�H< ���,s2����ڮב�����i���2C������%V���Up�o(u+�\��AS�T�<a��I��o����>�R%7�Η037ri]�z֤]�}��'j�b��D[[�I�v�,|,�����%����� {R�Z�k_��Z�(�m�S�rw<AV��é��5�!�7����쇈͗�O���	�~l�����1(�,�I�踄N!�a��3�l���LC�w��3ޞ�L����>�FB���;h�"�P���(5_@J�)�~/��z5T���l��P�T��rN�]f8X�T�*�������@��F��$���N�:���e�G�h�71��	�mц��dQjv�Z����|(͕qmm�L�s���F�Y�ť��(ٲ@���?��)��@@�[�qu�2�5B����R?11Y2WDNh�׆%<7}WI�s�9�8 Oz 8�����z�T�1F�t�o���ۓ���5��`�E9hэn��TS*w���a©�f@ُ����L��YZ��9$�`}���~=��'9h�l�8)A���K�a�"iL'�F���d���-LʚJ���*�jr�eKR�� PV�h�� =�G��{W�(�K]}&>�P���B��	�/���y�����GܙT��yf���W���YYH�Y5�ϚAI��1�t���C�KdfEC;�j~�.Z��q����-�j����z�χ�R�ޙ)�9�J�RJ2�
�I3��.�G��V+-{�;7��d��А�Yy�8��e�7H�9��MЍ�,q�6W�ď�)3�SE�s�)��^�(�������YuB�I^E��/&���/c$!ɇ�����d��	�2�F�����t����-�V�Aw����n�5O1����CV��Oa8�i+�sS��i�`C��J��,��9�V+��ߏO����^�����1�!ۣ)[#��<{S:�(�T˦�V��­��3a��|@U�Ip�u�
IR�&t��
���?+8���߷I��HQw�R1w�uT>��jF��B�c�,"�����t���)���\����*�d���whzA�f��=SK�[�Ȋ�bl�������@fw���P�2B4��aō�� �bgX�qs��z��9A�?u�q���vpj�]��(�?���?�}��5Ow<�0���$�nKڨB���o��'��M3��5ąQ�=�m���A$�"y�Yxּ�F�;�����
�ֺ�E�x���ѳ|⋨��E�ސ�ۋk�m&�r-�?�^�#�.��e��XƑ}�Za��;���9l���I�����!ڀ���7��"�P�=;�^�@w�'� ��	�oNue��A�d'tˊ�E灈��8�bҐ�2+�aY���%��4Q�{R�(�q��%�����V ���t��;�$zvrX�겉
�����%j���4��U�b��̇\Pԇ.��V���|y���h~����ß~���>Ll@)�����*�Ϝ��륦����5��p[��5F�Jl�8w*;?UU㱃�S��C,���ݐ���v�~,�W0�A?��?���#����Ko�6�11��@�֐:ٚKÿ�P1���g�#��<��^(r��W^��]A%X��㕹~�Q�2���p��o�Y�1��V7y�I��Sf�z�棲����8à�zr��v�d�)�Bq��.��k�_U�}�3�f0��L��Ƙ�9Jac�n��=�鵠�f���;&<Jn�<�?�QƋ�bY�P�Sv�u��`l���W�����-xPc�_������n8�1ţ,��FL�1ʛ6��ϏQ}Hv�`�.�d�����yj{�|���?�(���PҺcԂ�Zf�sj|q�
$�ov��M���,Aj�
���/ڌ)ء��z����T��d�x[楓� \m��B}o~;::�X�)�3b�<k0��'Y�6J*z����S䐑�yc�{-(���%��'�F����x<X��`>rXXy{�;��nK��<Ya�`�$���:�\DM?��g�n�aX��GK�STL]:�(��1%+��4�Ar�:BYr�*�U縮��Z�!����T��a�o�bY��r>(���T8	�~��ƃf݄
n3P��8�;�Ⱦ�7���>�.Nr���J�(�yX��g}�_8=�p��凕M�<枌��1��ﾳ�E`?�$ą�Am��I62�Ep��xUĊՐ[B>8�i�fW�+:��Y*�I�-[)�u���]����+�sV�,L���ʈ�5)���3�c'B�2l/�)2��L�����{1�͉m��/z��XW0S�#�����a��H�����#/<���d�ﳹK�$/nӵ/�/�ɡs?Z{��~���l���I��lQ����ME��(u q���)��������x=���ƍ��ڿU��FK(gЃ�Ҩ4�@�CW�x
���Y ��sA�*hP97����nmO=���D����_.��%Ξ�@w3��e�����Ǘ��kj��HQ�B� YR��ݬ�w��*���8�{]/��<��o��{?�0�/S0��m;�u�ѡ�c�!�2U� ��%�@�9XO~i5y���$ġ$b$��Iq16��X�"3W�s����5Y?���o�!�#`��`<�H��7 Z�]����%P{v�	���0_�(����$��ŧn��H)UQZ�}8���hᩍ�o��Q����`d���W;�=x��p�>Ԇfq�l�ڞq8*Ū˰cTf/�\�d�ad�	Ğ���,iI� ��.O�$9~GΟ@
X���N���hmǾ�u�� �����n2l
�`�Z�3��	 >b��m�����,���(�M%�qXZ�d.�J ��
��J���φ.���˷+N �:u�Y���_٭���+� �����Q"+��`���϶{���Ӆ�нy%�7��so��@h^]�ߕ��U��/��	A;�j������Bo{�=p�2�8i&q_�;�~%�b�F�y�~a&�ԯa#��5���;p��^�W��*м���(�F��A�L5)l��%�WPF�k�e7u+�UX�C�`*xX�b3���݋1��X�7���4���"�.��Kϑ�ъR+?*n�����)y��{hܪOvf�lf��0�*h���J"��P����(��MG!*]�Ҕ#�t��~��s��{�̓�{Fe�:V�&�� �~��!泵��*��ܛ�-�m�i� �J7���D�}}Dp��̀�LRήX��
<���*����d�:%s-��]����Σ�i��xӫe0P�W˙��h�Ѓ�����W4�y�x�	x��� #_�Dz��;>�T�g憭��.P��0)�kt�8@���f�!��D��]dss��Q��~�O :�+�XBI�@���v^Iw�s�C���CS(��W4Z:'#&j�����/��]���D�a���R��崤�80QZ�i��%������S�NΒ��n4�ɨ�L1�^A���gH :��a�r�Pד�h�Z�{iDdx5;����D ��2!9�z�Z�2Sq�$0��p^�\c�AC�z��������pP�Qv@��˚��#�Urw��%"��H'�H1?�z�^�='�*�syqz�Y�摟*���C`f��@B���7��ma��$f�:�xV��A �U�T�)�%!cm�-^fe�q�#�v��?�^�^��t�ȷH�S��-@s �B3�!��l��t�3ߝ�&�p/w8�����Ej�l�
8�G��1��CI��AB������@�3wR�Q4��V��t�\;g�������..�&i�r��½e�+9������sps���A��1���sr�U��+f`��D�Gg�w���}��ѓ��;�]��
�f\an���Qp��	I��N3S��=�ډ*O0u�0op����?�� ���Om������i����Q��#'/��n�#����ߙW�����ǈjP���<����?��������u�@hdf�yZ�P�lb�75%4�\G�A���NDK%Ϭa���:7���Nt	���$�ef'���T�XR@��j��)���D[ ߣ{}a,��*׃E�u�U�}Q��F�>�����OHР��{�sq�G�kR(��7���:��r�g��W}�aW��O	,$�!)�����x��4R�c #Z��5�(t8��ض��M��=K�Y���|�#7�`�8���F���R]�tS<�v9��N�C��Ҭbx�5u/S���r�o�{cm���� ��hL����i���CEʜ��+���t��y��[YXM�
*����������X=�����M�(���TH?x�$-N܉f<{P8��
˳{����vdEC8�����:�� u��?Ҏ���U�4�ę��z�h�g"�q�X�H��zL������I�<����Q�ɐ�G�����N����c�I�Q<������?�8\w1����t&��G�!����:V��0�PБ'"P�����-?i:A���� �W���	���� ?P�pD2�])]��D��g���1�L����y��B��K�Y�yO�.2r_��G���m+��K�S�47ֶ�	jz��FR��7��}햨^׷[	˚���58	t�R�ͧ*�
G|��<Ϥ���	���J��&�Y��~�nC7Y�B+��B��</��8j�O����NĿXT���r���"���<�Nx�,����Al�S�nS�;��b��R��բj!�_f���+>D��M`�^	�;�d��-�>�e=��6����E��jrU^}�w���X�J�&cf"axB�� 5
�4���B��h�;}{�Zw�abE>f�J^n&7�/r����A�K<g�ٮ0�F�݅�����gA_�K�)Ey-���I�VB,Mup��{��ƀ�y7 O��k` ^�}�Y���X�#8�[b\y��c�����NGX�d��tMۼ��ʌ�����+ B컆�&S���V���o�m�A�K�*s�c���F� �>U�2	���ay}L����!��;��ϧE�)T�!-pi�z�ā�X_�@��R)I]�U�(,����QpG��U3�?+9�����!��U�lq��|E ΙV��jMM'��T�6�{�@��
�(*�I�7�ܯ���p��g&�8	k��+�߽-Ux�����I���N�kG�'��]�nt4:�w��݀�5/�i�d����#�J1q����#2�<�q�+��W��.z��ʹ?c*�*�Vs�(�<�%%[�؝H^���I1�����}c����)F���ӱ����X�^�@)8b��Bh�(m���g�{=lf��ٰk���&��&��3�]k{�N��<�²�@
��fq歁�+�O �|�� �Ɵ�Iu�"�����k�k"6t������sCR��稉���,��J�<����p�_V�����]�z��ۄ]"dS��Ϲ�!C��=C>�Z�O��4�
bNGQ\c�~�/ �y���(��o����B��c��!��-oŅaܦ�G}��7�l���f:�a��5H#����|�xI~��h�e��H��8�����:�yH%��A�s�	�����Fd}�+��o���� 7T�o [�����J���Ƈɕ=�Z=�'T��!�/�*���qa<���#�C�Q�҃����o0V�)��u��ݡB5�נ��3�2V�}������f�^ ̥+���d��D�o�������U��B�z+���Gde�B|pP����ŒIpy)3��&Y�R{tm)�����ɧ�}�;����f2���/��X,g�Y�hx��(�� ��Xݼ�Lz'"M��J?�ї����Ž���ei�s�G���X�+x��6�_FO��4��t,,���Ft�W�����9��"_�n�Gҕ�X��6�%w!�"`�q:��/��|L�����$����3��Ո�J5_V��j�><T��h�DP�·�[���cP���ͷNe���8�x��(��m�h�b�`8���_Ɉ]UY傱\ʍ8���h?��܍f��&_��`��μ�Z�ܪ�ǈ�v���:���S���U[���(8\ ���q��u�JG���9?������5�y���Pz7��o�icNu�/�<�|1��)Ә���qn���㥧a� ���x�)�.�f�	\�(r2�($���kv����];_RO�CGi �5��N�"2Gڅ��m.u�g�E<������F*y,��l0��Y?�Od�v������{�s@i��9���䳅E(�4�ϥs�m���ك�%���3�
�fh�l�vn�aFG��>\����v����֘t��4�4wYa�x���'��P����x��m/��9+pK3G� ת����&��8�JpA6��KEIt�q�e��d�8M_�Y���;���aE}��G�
�o�mAN�a���;.�'��r5�c�[��{XF��MTRd���tzy��by�^���	����b�1<fєy(d|B���x#Җ�U��~�D�B+W6}ݼ�c��+-�Tf�$V�A��zMR)���5�)�Q��nC�\"1kĬ��v�wu�A�C���p�L�\'B��&Q���[���Y<������l]6���L2!��}vQ��Ɏ\�F�E�o���?m�]��ǁ_p��|H�0���Zh�c^��e.�a�[6����2A2���1θ�0����zyʢ�$
��ʋ�.���o�Ѩ#0N;'D�p���[Z�HXX�L��Zs��������6��QL�&�T��)�-�W9Zu�x\gBO�!���~�����f�=���� )v�x1}�����jp�%���:ﱁ�c*V�w��'�50�B��:��p�VD� q�l�\����.�S5�Q� �E�����ޢ��5�������pcIT��7ce4C�;.76`)��R���~-L]g�ph��:����]g��F��T���Oijj�3�(��:��)aIa���y�7'CB�yU�V%+�Xq?����	�4-���G�9�J��P��C��N�>�$MNm=7��� 򳾂���`:2��~�0y��L���;8�6U��V��Ym!�v���M�S)8X-*��X���J>����*c��s��G~9\��~lS,\F�"%ƺfJ���8���:�Hg��O]�q�2쒏�ct��e����#��7J�+�4f���=D+=.���M�B�?�3v[ӇȊ&~g���)@}�pP\uVV�X���?��ui�gڤ�x���,�>	�\�)��#E����3J/��b�G�6�8�[GT�aUgn�y��\��P[���lػs��i�\��{�^�a(�<£g>�փʣ���Ubf��l��ȅ�3PmD�x���O�{����y?�Ƥ?�rL����E�&��}��ո��k�LJ�	����n��	������)exB��FY��X+T�?q�ne�H/ }M=rp�K�:��V,��|��X���[�� 9���V8w�_=�1!W#�g�%1�D�gԵ������WfCn��piM�����Q�a���c�,q�bT`�wt����UJu8�9�+��8�L��ګ:��)u�y�y&o��V�@q�6]��'��y�q���7H��@#ZK�N�\�PL��v���F��P��u*�Q���
��$JA���g6؈��ى��
"˴�Q#�RnW�|#� ��4��||��(��*O��E-�(��'���B�@��q�siq��[���E�s��6����M�9� ��<��\�;�,�:�N�ES�F8��צ��~s����)m�9/����;�� O�s�aI2��}�i���nYF#$��|q�*K`�m�,f_f���m+�,�Ƨ��Y,�M$Sź�Y�>:�tۚ�y1��K�Ϸ.�p��2�DZ'� ��6��|��}�����'�@D���C��.�3�����*�B^��(|�ŉK�OK ^���<�6�lȋz=M���"����I^aD�E?y�W�/2ݮ�(YZ�c����DA�� #�C�A�G�2<�Ŭ� p��V����}`�G�fg4��ψ�I(���9ʜI߉�I8�����ag%ZkK�q՚��>���}�8A#@Մ�X���v���"I�#%�������fU?�yN�������W�.�Wt��z�lՋ��
��<:��E��Y�Z��)���%|�$oA�v WI)in�-���u��F�z��#{mպ��|�Z�l
�0�������-�,������p���y������;�k����#�[Br_�� �@��R���\(
��U+�k?J��o#��s��9�Ȭ�7���f��%E^���d�>�$[���F��!�銱�<����]��U7���Ǉ�G?b`}(�UI@ޟ��Ң��x<Ob���`�]c�9:c9P��I
jd�z�
AQI~D&�����e�]��K����uC�p���\��Q
��|3_�s��W�$ɕ_�E�L�@���Y��\�˧��f���]���	d���� nVl�'��8��f���R)��61(9��_`8��
&v��Ԣ�ɓ���Ƽ!�����Փ-�0%�ڣ�iS��4�A�"ض���N�k�>�������ہ��gU���EC�N٫��)�a׮c���g�tIi���EW�#^3��0|Ҿz�w�<��M���Q
��"&~�E��Q����Py�E]��%J(�`#:��1�<pU?�ih;1���=��Oν�2������B���4"4W}�`���@DK�$�n,k���c�^�Y�H��)��:F�;��
-Y&�����l��6�c�V�Q���(��z/^�������сJ�2�{(U2.*
]�]�.�!�|? ͕@��m�0�����ox��~�-����ݸ��wm�31�y�"�{���"�TPR�K�/8��C�s6�h��v=���G{j�RH��e۵H��:ԬA	}>�M��R2�W,�SR�����g��m�rq�h��T�j�?cm��5�&�>v�6���DQU�h6��,J��pY��>��A�����[[NJ���F��-� ް��C*1��p:S>��
�R���rg��1K�B�VV�a��a��B�j��+�ǆ��kt=2�>^�%��S:ʮp�<�H�aFa9��1[N,� 1�uw��55�W���&��Ͻ�AV�xWL|��y�dkNKwy
�ǃ�+�L��@�q&�3F����ձ)���\���m��KwJ��_��7�.]�M���~<*��"��{t�$sǾk;q���Fg?�n�l����1�p����V+Z�"����Ml�`\���;��Y(�==,3�e䯝j����.����|��|��cG91�s�0!�\2_��-ܱͨjD�p�gk0�A�:�:� �,�P�E}v�f�^IG"'֛���2��<�6�6�s�jZ���I���z]d�f(��)d��cIn*����F�Em�J��]0�0��������OU8.��ոs��v�S
~��~�_����wC�ql	~�R��'���#O@ڟ��
VS[��#�}#���&ɓJ��(:�����
6�����*�w�,s5��r�L���������C�feς!�c[-ş
;tO���"���1�if{��u%gs�vl��O��g(��ٽ�k\H��i �����Z��	�O��u|ډ������ھ�Z����D�8�i�_������v�]�74��'S@;�����xOZ����`��12nF��5C��z'۽��%�Y�^�\ˤ��N��*�춅v�@$X�G��X!���hkp�n��!= ùi����^��\ʍ��z��t��^��F!3m�ņf:�;}@n�ͺ��р�|ÙG���1q��$�.��`xy����:�m3]��r]��>�`�gخr�����_"g1�g^ӭQ��]�b8���Ga��t�!�����1/�L[�v�y~�
��D�?�y�@
2���q����7��v3m�*��C~�]�%���~������l��4b�p:'L��!Qh���w�(�6J��T��5̓qX�F¡�ɫ�㐭��(�|t��>����ȓ,�[�EZl�b��Zı���Z��M5�J����	�r �Sdj$���[�.%�I�B��2Spx
HFױʩ*��'�����`������8�`��e��|hM�G�{y0�b�v�^jh9]�WK�����d܏���RB����;U1����N��|�+-��W;h��V�@=�)j�j;@�#,C�S�5jT�ߍD7O�މ�s�ή�����9s�!�֖v�}���;���b{���U?���[WV�-��<�t/W6��x��S8�{f���7�uo�_������>�[��Q�~�:�}�͒0�t����a[�,0�JG�4Ob�rd�H�x�m���g�K�"��B�g��Ǘ������?h-��h��I�"�A�(�LIV�HT5�������!��C��L�ubk7�,���q}��8��A�����0��k���֓Ի;�;�m|/����<��F�ƴ r�9�m��_�N�I�e(܁H��|����t�	�s�ɾ�/2�^��������C_��,eI���eNN۾Y �fR�J'��p�}z�~dqg6<>����X�2���5!^�Iʿ�O�d�:[-gK����ݜ��D?T#��E�k_�9��g��S��@�Q��X3!�i\'�=����j28�4�HB<�_̠r�!a���O�n���C�uJ#�k�}(��	?�k������r���{�T8R:@*��,"�n�z�]z��QX���/���#s����ܸ�al��$0@kڱi��� ���p'�£X�Oҭ�6?�VX�i����T)��_���Z� �X������n��P���8�� f�I�:+P/CB�g��M�P��o�S�A׉-g�?��[ԊT��DY�.�ʡ�������Ǘ���+��X]����Ir����VdCCKȓo���8A���8{r�%��*)��6�����Uֆ�6�L�fJ�	Y�gL�!ժ1�Ϣ1�B�Q;f<_w7/��b�q����h�Ϭ�[B}�	��DLW��@����z������Af�&{A��'ai�f�Lb�&��	#q�26U�zQ�����$,5��q<������G������a��\�Lۛ�E&P�����"��!욳�5�g$G=�^E�����m7'�X��*���Z�	x�B5�kaj����yW�����lpէf!���.�Pft�	�
>S���	���WU+�OO��Z*8>����7a�=KBY�5�+O\	�y��]3'��=P[��>�hD��G�?��K�k������کx�t�B��O���L MmGBx�1�5�#�{�t|��.���P�S(E���E�ns�v5[�$��ej���cb0�XdhT�������=%K�*�O��	��~OT\N�0A읽(!�$
�Q<'�cf��ߛ�� $���Hp�=�ף&1~]U{Rj*�ܱ�J\9���#��|�����;�����D%Fl�](�����������@X7�/��py� �h��6��P��^�a���}L��mk�඀m�U�10��5,PF��+�>��/�	r����R��)Ιt�?�	��Jd�����>?���q\�v�D����I=݀Q������㐌s�c�[	��P}�љ��0��'����[
���ڥ/ ��+�t$o�t�!ώ}��,ꜚ�MI�Q,XPd��A�S��u�x�D��&�@4��1{�|��Za눥���KTa�Oє9��J�Tn<t�j+�d���qI��}�\b���I+Y"�uO�U�q�餥�s���t�N�g�T���X|�x]���iDԠ��s/��������5q�i��^�U��8���}L�+��� �B��6jy�籫a_K"+s�B&����b��|����=���E��LNU����M�3���N�@�9�����-ji��%x����ytj
�H�T~�حPr�Cp?gm�4�\��D��2-�3�.�Y�h�L�[A�"�:T��4B��_��蹏�ռ�>�K���.��c�x�����Imwa:Z;�|)7�dK�������b��B���5J���|n����=�i̟s�h�$�%I����=&��4uʳ�xJQ�Ƹ&:��3\�UPQ
�^��/���:����
�{����}O�[��Ef�����[3���[����{�t��97�a������:uԕ�s��q���bYzo��Ǜ>�7q�߹8x���߯V�.|��x�*�>��M��c���:�f/*oB� �n{Ҍ�C�{��`%3����JmH/O(��W"����kc����)�k�)a/ңZ�'k�
C�+@�ъ�J7K�ra9�>ՀI<��"RT����*:@�{pYQK�{�wD�!�$����T�ɜ#Og(4�3;g|�Hc ��.�`����-�����_U
 t�h�ɀ��}*��BzJ~-�7�P�i��A4���P,5ڲ�j��.W���6�OjD��(�3��=�-$�#/��"q�T`[#���53����Foĭ�ц	��*j���w�]���+�5e�4S�Dhкm��3*��n|��Rd�U1����^�q����G�z�]���`��@���{�>��0|�B�o���ͷίc7ق�}���-����|�g?��%`¼���vhDLS,M��d��'������d�*��qm��W(}������IĐ8ey�X�@��껥|C�U�jǝ�̋����al��֜��i��̩�����w63e%��p^q���_�P�~�����@���ϬQ�������*� �E\��������-��h!Ѳ8��[�<��;�#�hJ�������[���si��}���2���-����?��a�&��;u�@���H�-o/�U��/��%��R�s�P� lB%FE���1ܢ�3�J�px~1���L�����(>n�+ƪ<%8�����D	,@�(�
�%Uݎ����6�/��~����#�&X����-Z����@[�A�|嘃�?�ĚӖ����,qy��uq�M��I\�\ϡޫ�b{�ow-?�f.���o̡�z�P�=z�ƛ$��
^�T[%�n�ya��'U�!0`��t1�]��J�~�zK��3��m�A8>~Y5�1��O��e9�	i�z�]����"c������"�E.{��&b0T��8j�S��/���=��SdJÓP�����BEbs�Zb�1���%�xn�V��4�Y��^���Ym�]�j��E3��Ǔ���E�e1�Pd�+N�k�
��"3����uaK	}���5t�
��A;*�i}K�}��K	�YG.\%rN>ǡrPs�#R˰�n�Y�"&�F�{'�C/}��K�r}�x�`��,�G��?�h�pӆ .��� �.���d� �s�{xx�
i��EtB�\��Q���0qy/	�n�`��{�=5��4~��W��<�}��������|T�о;- |_�m��� HNM��!���iw �0����Jc�m/�^Z���jzT9��e�vԞ�).��R�D�,`u�lK��}� F(�%���W؉��yl���S%�{�B��s��k�s��6Z����=^��/TzG�*3Ѝ��o^��u�O\�9���EG%-h��q���{�$��5t��u�+��O�Vs��͋�Pel�QԖK���[���ơF1� �SC	���}���u��Ĵ��������y�Ł�VNE�GA��غ�a;��:��B�K[6rTݠ��2�j���op]�_\��$ g�����h�����o�|�3�Ͳ����=;9��b�������onL��E���7Ii=��t�YD��<���k�C7��v�:��ʁ�z����ǿ�Uς�7�?%������7��3���l���H`>� 0f{��F�my�t�����Y
���1l/�Ŏ����``3��2��Z �4�q,�)K��K����Ǳ��-��V�K.�~N^#�č�e��4��T�����ufuY����~b,:`�/y{�R�C΍�X�زfW��d��~���M���!��9.��e�I:��}D|��R�O��;�D�ҬgWW���5��:g����ЮTeQ���XHk�yO��8��]�����춮�?wj�����0X!SQ�Ӛd����!�K�:Ə@��v	Y<�^4m��s�
��z-^M-��y���g6�N�`�|H��,��a~�n�.���c��dݶ�"�]��N�^х���f)�g�P];�%��O\������^��䳹铫�͌�1#�b�rQ�����cp�
��K�]�d��#�}�>�o��k\�.Z7so��`�>z\����+?�ޘ8��]�<����!�h%VH�/I%�<h�t��1&DFb,ʈSS*��� �"�l6��$�P!��*!�8����Y���}�G<4+�X��m\�ٿo����H<���= B+���}s�`�N�n��-��ھ77K%��}A�W�jӲ4d6̺��xC�T��wB�%6��LQ��.9��5Ї�-��Mr���֪�ߵ,����"��}�9�kz0�w'3�t"�0�O���;�jɅ��� |�Jh�t��9$�ca2�u�����h�:�K��	�p�a��A3c�9�M�x��ɖ�/�`�����4
&*M��Y��rR&�YӺ@bZ��kUa�/1Xg��iU�+����lM;�m��ֻ��� F��=C~l=|�R���VB�rcͱ�o����|x8,����	RHe�)@c۪$Zz����[n�f���J4p]W���!P�@�����1�6 {�*��y^:�&/U��&G�a����P�p�r��y�a�^U�ZI
�P�q@�'=�RR�dy���*��n��?�V�||��y�ԧ�ؤ�������L���/����t.$�epjB_b�� QH��%J�ބ��.cG��f�eѠ%�:nρ9���٠0�g���>3�}��<|���wS|�����kA�W��q���_�$��I��@E���e��:�]'HLmk-�ߞ�g���9��=�e��̀>��:G�l\N��g�w�͹�i��{��d�5NCB�c��~"�>G�D�� S�Ψ�<��ʨ̸o`��Z��k�� �������bdud^�Ul���[$�q[�{y�wt��X~���9�dX� ���3O���18s���rϻ��z[�y|��+p#7Rr�~<e���B͈i��Q�G>,�83�^R��5��I��G?`r��@G	�<���SO����	�gGd��&I��8�p��'a��b��3�κ�*D��;����/|Qʟ�{�:�0D�^�dy@���и��%�Sw�ƴ+Ŭ�\ "����Jc����P�H�"RW������o8S�m��Y�t�Z����Օ���6��"Hy�ؓkY��I%��T����!*wZŌ?�i�KG�ΐ5uBep쿎X+�\V�|v�MdX��ٛT���'�n̲s��S���Ľmqg��%(R��^��:�ӟVH�8�k��c�=8{G���($��]�C�Aq)\k�G��F�Ds�+f���z�2��r��R�k��	��ZD��C!G @���b�
�L�0�.|�~0*/fh��HQ��{��Λ�h,��D{�ac�OJ�22����`*]�s�ӎ3VF�@�����ޟz��w�ĺ�ip��:�a��?=%Hj����S8i�hS�����!�IC	�`n�Ͳ�������%���o�6�B���L��E�1@�����#��
�޲]er�_F�%7����w ,ZkS�	tP���`O��kBȺ��	kRv��ჩ��*�B��%��e��k"7��Wg���)��E�9�*ώ�H�}���"4�����0�%a�sy�A=up�ȿ��,+��<�j���mm���'�����Sx��;ה���f����U r�����{D�	������0=�7w��"�&�u��5�����憾]N�kR&5�tt�дw��⢧|�6����d�W;΢G�t��Q;mi�y��T�oQ%{��p�������ۯ�+W	���y\�P�M��\-~��S�
Q����WCI�[?ƂO�S+P�L���+p��X����^�9J�Jw����~�+��%|;��G��5Y�J�%{ߏ��~���8QxL#Ohj#��1��D���.��V`��S��/��U���)��a�w���%�.�D#��xA��IcG���ŅT�_�|�+'����m�H�E������Zw,�ǚw>��Ő�	;�GZ4�.a�<r:����:俋17١���D����7	�98��Y�a|���E�
��z%�{dB(�=i���}��.�Dg8����͢[Z�_^�.��c��6�V`=�H옮,�O�$Ov^��
9�\Yדڴ�o�I�]TS.��ܴ'�f�u�t$��M\�1��P~�V�cuN�lz��/_7��ӊ�� �5OA�� m�L���Zx���dY�,~�y�{�9�m���V�3�w%�j�?�:Ϋ��\o!o�ZRW�p��?����B��?���=�68 �T��aT?���0�~�e���#��7��ٰ�*J�#Z����A�m@6���/[Q�9������0x돛ggV�d��QX�p������p��p��:
���餙�,J���n�AZ��.�S��re9�iqF��9DV�µ�-�׶)�+��E�}�<�5�J9x�{�u��e	��\`��.h
��4�)�S�O����(	qy�� ���2�I��v�Iڭh�$y��>B��å��|�jA��^���t��چ���Mu�eY��c��֙�b��=[<g���8�j۷a&�Rf��� ^��7d�#yt����C}�~���gѩ�웍x
�+m�#��,�ͷ��v�'˙�0�n�"$�/�|�&�rsX�Rڃ!"��j�� �p����hx�.���I���o+\����{�	}~{����(O2z���$uک�)�X/R�D+���B����9w��1�����\b5u����vwş����&�*�OBsZ<+�%0�ٞ�Dns�O�:�6�*�c,@�hmy)���r�"^�@a��k�$r����kh �s�l��\��M�Pݥ_'�j���p�.饨�<����,���;U����dQn9�6�-#O���Z��k������G_�7{�d�¶�;޽��rw�Z����D�G?r�'���$ta���7z�N�ԛQ���mx������X�K����&8��]�gD8i�w�5�=�D���T�;���0�ˌ�������{�PeE�\��_�J*�J`�d��"�4���ۜ��?����ǁ�k���)|�I��zK�L�-�N��������.2�M^p`����հ��J*~EZ��N&U�j��#�q�H��߮6e>[ l74��zsT-ćA/�`1~�	@z	(�*�qq��
;�H9}є��(q!0��|���t�˪I�y#C���G��T&g���_M�0G8��禃�!Jӭ���՗?�&�zt�Z����Hk�h~;>�M��=�,��:����Xs p���o��Z�U�ߴ���N�+`$�k��ӡ���+�	h�H����U�V�#����
Rm/AdX��"�F�jG��Y������RF��sq~�]?ܤ��p`�����g�`Z��`%_
�:��J��n;�
$Ƽ�*���C��;���oQ�D(��9���=�^�D��c?�E��3����ʮ��g����!B'[������_�&������,�����A".�G�ԝ��FP��L�3u̺#O�����E�$��B�&����f��(GZsƒ-sf���+�Nl�A�s�m$�m#�>!��xlX}���h�pڞ�^��W��yQImkA�Ӥ8����R<�-"�3�/_���L�./8�R��尹#h�{9_FА�R��ɬ��¯_@��/��s2�(N�z��c��#�F������)n����F+��F�#!T�bk{��� �ι9��λ�_��f�M{w,����beL��Q��?��dL��a��X�+�C�v�v�vGwt
��B��v�JcN������j���Jܐ1d��Wg_��rt��+c0A�p�e�����'K^��c�j�Ax�3��sT�H=�2��$�H�D�@v���	���U]R�	�H��v�'���o^.�F���}�%�j�!I4��P<�0՜�z��R{��ׂݝ�H:
wC��*�v�[zv��
k��6b_B(հ^���[k2h�D��W,!�tO�+�M�3�(.��i�ZT:QiB�~�U4����75vM	<�S5!���)�Gѩ� ���ˀ#���Y���;�AK�m1��q%E��L'>s�X�>`/�l����	�j�Bfs��e4+�3K�����oO^�<�!�����(�
�l\�T⍭P,+È/\��Z�T��YS[�b��m���b7鍹�NMW��j���O�	<����j��2ّ�Kn�Uuԅ/�3�	�����Tc] D7I,L�bʢ����5���%"Y�a������F�Bc�s%��V�:�B���wz�D�������_�����X)�Z�5�k�ﶢ�)QR�1�DD��R!
�K���
dڨZl�7�8|w"��X��}���E¸�N���ڨ��~��ΉQh1�_,�HG�b�C۽�?��j�������c�$�����F���'�د,�֐;5�b�<Z�1A؝����߈bL�r�\�S�'d��a��ְ-F��rI��۵��.m�	t�%Ti�y�l$�I>����/�<\s7h�y�^e�@��>n������C�aX1@�/?��9I\ΰy���2dVc�a���;-�~���i~�7��Tz��,����e܎{���-Erh��0�f:�!���/*}��9�d��K`d�^�PMV_��j�f]�g��θߖ
��Q.hm�+��O:�F"�b�7�����b����ɦ���lJ�^�e�|�USP�������0{z�����u���!�&�ug20H_�;���vɒ���{ �Ñ"/�Cʛ��~�~���1��(ҿ�
�Z_�Y\���ۄ��6<`#]��)��܎�GID<IJOAa#�����idJX��=,��p�uw��^X)K<�6�z~)
�M6�y��Z�!�'"@/b���`3B����r��M?#,�|�`Q.�*�
�Ho�,ۢ�h�Xf�i�
t�QZ����#MDI�wse�+�c���<�^u�� 1D�][I�e-1��� ]�ְ�H�����ӵ)W �Y)�ˀ8�0��vl�G�s��`�eqpu̒�z�*��Ff�|�9:�A��Pݙ���-�Cn�j������I����&�����\L��(ǽx��p�-�RX��vX��m���a�|�B;�f8�~8:6���rI	ݟž��6R=*8l�_	�y�"ʆ�Y�4���Ŵ�d$�C�*�Ǧ$i�N�V�6��gq�P��LO�������\' �T�_��cm8�����=��ܚ)�?#��=�F��`�`(�~���ά�j,�r���R��m|n�*N �`�u����Վ��|_=��z��ͣ\�aW����'u>�~�%Q�a���tY���RP��8�P�;'u���⟉�l��umJ�.����0T�`wt!��W��P��A��K:w�~E���`��y5~3q�r� ���>� i���Ԭy_��5Ɨ&����?��2.D�߆"�bR�9������BZ�*~�y7J��.��+�U,��
�q�r�PED6r	�B~D��U�ŋeԧ8��`�)lϓ2��n(�iԒd�>�e�D^��}.+"���K	��̐�r���v��^'p����l�y��Z�N�����ƥ0w:0F~�y�xߝ=�i�E�kPbP�W�I�r` �y�
V'b+9���^F�{�+}������#�Í2�[?�3��`oE�7�""Z�ks�QiY$��vV�E�����VGO��� �L�'�ćw��V�L�u61���@0d�qHTӘ��� oce9Ĝp�8z���� ϶ ���^�)C����U�Q�<��6������N�}��f��Ӆefr��;W��a���۝.�	�o%�P���ʌ�����9[I2�8}�e��:�%Y8�b��
�7+j�^RTa ��M���q����D�E"�޺��7q΍��̣x<�$��Ofs�(�G�vݖ�|��d��\���<��}tU,��n�j���6p�<՚��q��p+{+a,#�yD�0�}R�!��#�b����X90�7g�3%=���ۓ��5�����=�r�*�P��s�ș���D��d,�5@Gq{n7�%3�C�%'��.���Z��k�����%�@�=��p���[��_��y,�OB:av�������?��u�z&	ʠ�K}���6&߂�9��Il��1F�S�ml��P�_J��^BQ�!�����}�0|#\nOyecnt3�迤���_G`����yt��L��Y-P��VҺ٪?\aR�+6>.�k�,2�|R\L�2��k����<V�#�=ێ�B�ϣK��ˮ��+����)�jMf�W���SUZ2	4���$ܒ�۫���w���^�|���Y6먍8]?���~>��6�t��$���X:�u�(����b0���ɰ鹨�EW��>]ӰH%���q3nBn�c�Y��[�g�<��Ƹ��v�ם�X�L� 1:��֔���=>����Ĭ������(p�
V��x�n&��Ε򆇑�wݶm ����7�)9�8�L)�z`H���] ���y��3�W��Pk�*����?��x�0��͆#��e�]��ʊ�2.���`mS�~�A���UoM�-�pf�p����yO�<ە��s���r��Tg���jq!9��ko�B}�R|q�_Hh�m.�͡��*��"��I�p�2�ƹ���lۓoq�񝾍*���$�~\)�4(T)����iͦE�X^}��C�|�U�(n}��EEY�C���@�h�R��.Ȯ�
�w����6H��i]��oD����ho}�XY�=x��1t��.O�\KH��Y4kS��=sNf��Ja�/[&���T�� ��5t��>���j�����9
�����k�J�.d���ޯT���!w0�"|c�k.�G�����$�[�CHQ�V�d#�V��C�����u�Z�YV��
�����F����s���s�G'ƅ�N�B�l\���˂*�<��5�#	�E�����kT� ?zfZ �˶x�����/�bQG�4�_AsfF"5D(
:���:�0C���ޞ�|��
Io���d��͂v�52�p�%�H���@�Af�
Ö��]��������JR�U}���m.��9��+�qO�h�'��pʍ�i\�#�� ���-w�L� �+3(I�5�xe_o�37�Z&�R\h�~�+In���Q�S[���`U.f�]�2� $Sg��'�ɵ^�g1��48��W�.7Ȣr�p�R��������JF�}�����Ex&��$ :�5���vUD:�$��f�&�t���y�z9��a12��A��3�L�>s�uSt�dL�=�rϔ�.c!����X�z�R�����?�V��7>�OS�=}��ĸ�-�"�Ȕ����RlcU���X�m��H��E�S}��n$�D�+�
� /��-��.1����(> � �͌�ˆ�����q�yߋ�Y��q�f!�����%�eK�([		�c�09��"��hScd�SspR�f\�\͉Z.�P�{�iYb�m�W����=��8�e"o
�5ܤVwRT�e�.�M1�rѢ�H�Ī�����_zs`УȠ����>�F����(t�]m<���Eo'���Q6�$���[O6�#�������܋���[<C֠�Ԋa��p&_�o%}�5�C-o,=7���$=� ���<���'X3M�?���1ҝv@a^8�/K,����z���,����8�rZy ^�f���{Y�+�v��������A����0�^�	�[�_7��{|��������ظ�.^EZ�Xgsk_=�v��ʳH��=z�652�#�a�-u>8|�记�3�=��	�fD\��NоMC>�2פ.�:�v �d:5y_�d�N�'/��
�����@\�M2��1p<�h2�Yϴ��D�J��"�_N���ƇT
E�np���5�ͷv�3���َ�ȲG8���a�����l��	�O�8�>��u����X�ωg^� S+�p�gE`�>h�?�vX��Tٗ;[�i�_;��L+�(�i��8�@r."����hb�N�Yq$���H�@�T���g��3U�(��$����?Hu;!���^�I^N/{}�_�j�8O����	��8�"
���e�u��X"0H�"�}M�r�Y��OvUq��a��������������; �HӇ������+Q�^U�!��n�����.��"z��(X~�_c�����B�ޓc��V�|́�vft�F(@}p���wQ��5{�W<ٹ�P.�/��c�I��o���/�p��`�LZ��/w#{J��8���r��ĸ�2�=���~����EC��kgm� i�WN����7��G������ߍ gp��R뵿�����~<��$&�tG51OH���
A�PYݥ����N�G��R�"�:�`��D��4b\��u�T�9%��t�Wa�Ǫ�{*���^��ˆ~�Y����酢�b� Zx��*��x\V'+*y^��v1��z��J�e�K�{6�}�`�sߔ@KA~����{����X>r^{������f�8�V�/vuR���&��\��4�F�+��q��\z��x�<�8Y��o�����]��="�̌L0K���0C_oz^ z��g �+��K}�ױ+RI���E�t���#3��1g��Q����'�B �aez��l�{��b�u�@˘#�7%���OIhR#\�N0�����k�r��C]P���hc"�	���ܻƏa�Q����q%9�)�H���` ��z��݇^�w�o�����P��8��|,%qUq��m�4d$��6��Ѫc�,L#�f��bk���(�&{�Jǝ���P�aװY�
`�1.TpO���HxSk3�sZ�O\h �9�A�Ț�j%Qv�7�1��o^��P,��]�Ck�|�D�젡N_c��C�m�E߼�}����;�>���TQ'�{�=r��R��8��S�@r���1�Z��='��\��L)�A�@�L��.ak��B���GAz��K�3��PX�oډ�� eZЫ�}�ÿ��v͈���x%I�����N�V�[!>:ῆ��Fms�?M�Arp'bn2�/����fm@Q�F��#�p*b��a���</�3�k�/i�Kh��B����y)vL���&�4]�Ez�wO?�l\��O�r�����g�B�1 �VN��YEzv����7�"Zg=dť)7D�B�(��2���[�g��B����� �[p�O��ZsΉ:�74�ـ@�bxޙF�Q�}J<I('�!�깞�3����ˌ=�������qc�k�&?�%����uL�R��i3P�
I�e��ů��0�Vp�S���������JEc�x����q#H㊌<�GfV����\���@��t\_�G�v���A!�dj�v��CD�͒����C�@�v�����ҲM\���D��r�|��Z3�Mx�yf�]���j�ӈ7�{�팤���-_�r\
�&m���3�f3�f�G�zද�p`TM39�V ^��IQ���@�ݓ��g�;=��&kr�%��F�HCK��*h��5���:�8�Z�:p�Za��R��X����Cb*\��
��9�{�˥恢��kI=v���f4N�3Y_Ȯ-Y�y�� c҄�<5����9XB*�o��بEJ-h�K�ѳ�̷b%;4�Z�I���$��Y�W�(e "sl	�tM�R�v�W�#Vz���[ΰ����~����"~��sb��H0�|�D&�V��}B����[��{W[Yͨ،���ԴZ1����T��.�$��¾�T�\�@I#�0�X�>��ϊX��(dT5��|q���ReЊ�&mܦh�c��J��O�Ym b��p��d�d��1xy��5���.��&W[;:��Q����m@���X�ԯmI:P�휋��+�G�C���:�.���B��[�c�.����f�=� �k�8~/��p�l��>���ea.�w�lzVA�E7|�B�z�\�5w�[�&0Qq#q������w8o����_�RTMEB ~,m�̃SC��л�wE O����n�=�惺ե�T?t��±�4�v���Skֽ4��&Hj_x�Q�-��ci��7HD��.+1�кZ������d��Ɣ��Vv]|�(����NU��J�s��.�>870j�&+gl��G@��;~��[�p�"H<E)K���[�@<��zT��8w�1"�Y��'l�8��W�����jy+0$eb:ݫ�Ϣ��9t�;J" K�ᤁLɐ+d5T(]HB�	�ID�sñX�m{��Qt��A����*��
��6������q�3E�l?f:��5�>	v�̿t%E�`� ^ƌo���9�����$��y4Vh:�H\-�@}d�D$�H�)S���b�+_��ePi��f6�°pe�3Ïr�A%X�M��D�6$h�(X��5�U�j���}������
�(LJ��͠��p�$�}�z�Zi��7��~QM��8�w5��>��pyͤro�E3�tf�5��� �,�a���B�`��$��?�xܼ�yS6�{5,�ugrc��q13�z-5���+�Tw��mv��XI ����c�������Q-�b�wh��[���l�%��S�� �v"E!�
����͊SG:����.��o�s(W3[�k�!�E�T�{Gy:v�7�(�W
�)����4�/���W	
�˳�5�w���[��Zѓ��z��+�n)���[ ��Ys_�	Q�z�/�P��\�oK�\@���]R_P���gQB�$T� ?���X��u=��V�= N���`��@ת����Y�OH��^�d�HƎ��D/M����zo^)�U���:w��
yGⴅAr��~!A�����V!&x�V~3�����w���{�Ac�������_̉Ǒ4� ��x�o�R3�ݴ��/aYQ�9BoL�D���)�w�f��i�0�ML�Η;�!g�q�i�U�'�^s.����ӚWSpٵ�W���d��E\��I�O��D�sƾ0��6�Gj1?�����9�5z���i1x6�.���D��U7�#�ohbP,r��9�J��ȻS$�<rM�T�&&�R�ĸn�Zk���Q��Ƣ���I��cSX���Z)yUf��bR�`�_�	�?�m��K�^���ʲ�p�4�ϫa��w8'��w��Zࠖ���f�l�w�����mx"(�Y��(JhI���?K����|U0��|Ӯi ^Be���3�As6�=�+_ ̭
W�����>�Y�̬��	�.ޱ���ޱ&���`@Ȗ��J�*YGI���� U]��1,*�p��S�n4=n����Ǎ~���H��˃06�B���"$݉��=�Z��ءEnH ��t�]:�rMV�G�>�B)�t�?*f�����B֮ G���1'�uT~���4�e��Z'��gE�=�zD�Dǚ����l=c)�Zt]�1&A��^|�h�g���*P��T>�[��y�ꃡ#���yl֛wUփʗ���SvӨX{+�u�TNi�^ZoM�Nc+k���BJ:.qz�Rk�7pt����G~'�i^��U�A_$� A�P�0�	a��՗�#dQ��豬��H��U�����o,����f&	����!w�/q
�}s���/f{�Ww��ġ"����s�%�Er�ި�u,N�V>e��f%Mf%���7��6��$��խaa�Ns�د���/p��"�)�g����jK�Z<�(�Z!N$���R�vݘ	���3~m@/���3��fj����ϩ� ���^_�1W�����^�uɚ�?/g�T3N��K�ѫP�P%��M����m�xCkMΛ���i+�DO1�&
��`B��Q˦��<��(�'��>X�I�.�I��i�g��v�J���[�zp!lx�>�L�UV�չ/T%���+zWj,�R��E�ÓS�ۖƯv����|d���ut1��:�c�k��c��ɄO:E���_N̊+�8c�1q}C�^C��Q�O�����p�cQ;=rRq�<��07 ȓ�l�Ϡeㆂ�9߇�!EM~�m��H��C�2h�&1X.��m��Ǣl`rE�M������ټa]%���h�2]��N Oۃb�Hg�+6�xC�bF����!L��]�ttr�?�;� q�RѠ�F�i��]�<�p��a�`��e
��d���/hP����a�5I ����J�*l���*�ip#�>k���F�`��8�i9�Ң�<�Ry��r&��H���7��@�?�jphn�l����}�����9��^��Ү{�mm}g|ZT�����	B����"��]i�w	-�o�B
��n�{�V���/ E90�����?q�.�pB��]�f��}qr��F`�_@P��%׍z��}�+7���b"f�W� N��ٲ�s>`�Z���hF!�k4T��g/��&nn(�����݌,*����v�"�� �F��2��Iȋyб�ϖ�q�W��=�'��;�E�܅pFO'�����I�ۊ<��i�&9)���oe�K����_�/�&.R���F}o
���Ga� I>w�o�T@��\Õ`�s�*�{�Ƭ�����S� �>m��'�dzy��g��b���.�e"����8�[:
-;����U���
XD�X��N���U�b�Mt�"���,�#�x��1���*5����R5��f����~����Bٗ[�2O�S����MMh���X���=��0-�0�BkL
�0�aygil���|�&�3���WʊuB&d�O����"neW�Į��w�`<���)�<���y|?ߡ:��t"����~xp��g=��v��{UN\��+�vFΞ{ʉQ*C��c�Ą� i�'OA1T���O4��eK�m:݂�;k^��y�k�^����^������8�b��~��r �o*�V�j`0!'�	�]\E=�r�!m6[.>�U�_G���8�oVW�&(kMDC7��5��P���B��\�Q�C\�g͖��}�3dR�6���S�,�4?��.�}d��&~�k�!+Ԙ�e�y<��%�����`��7���>��3abKf4�}����#z�[{z��yQ=�z�͔P��oF�7hS�&��]j����L;ٻ)Pg$�̚&
����	=��F���kٜ�P����yV����\��� X��L�.�uu��n���K�Ax������pR�|�������,��Ut��5J�����r����,�[��	�=o�C��ᅿw-�p�������<'Yp�1$��|-Q������'?d��k2��tL�k�*?D��n	��L3i� �j/Iߗ}˥�!/qW�QO4���P�2��/�0z�����,���7��|5��Y�+�("C$kS�s�x��~^�!,��s���}ǴN�_�WbE`��+��S�&_@����_�]�����Y7<1�$�	��!
>��r 1wy"^���/�|&6q�ցP���7~�p���_���%�4���z�j�퍫<d�g6a��S�wLi���L_#���>�7y{-^��2T|8�DN�xC��o*w(C�c�R�$f��4N��r�%?���;Xլ�����E�'o+�[Z%��!��#�KDۍ��%�l���Z�e9��ޛ|A�U3���D�Id:�/u9gȣ2��ܹt�o����p^��1	/����n��p�@�z�����r�KoP�YA>�I��҄��\�#@�D6	�SI�����Cj]��5�I=j������.��$rSo��颟�% ~���ư����V���i�WFAy��ؾ�a9��('+_�#O�ɇ<��~.)���;��	[�p|��tȼ3f]��ٗ�}��<����#�H�t�0R�;�ެ`^
wH����l��/��h�#�Ƨ#�^ƣ?rW��o_���FkD.mcW_\f�5i��y��2�l������{^G�|��
��(忭:��(���� k�����t2�%?�t#<�%X�98���c=]ވ��o{�Ht��e�@�~��-8{+�NZh�����g%|i>+��v����#`�^7V��H�k�S���	�%m,L'}��Y��A��WX��l��O�M�x'��)�%��1/1ҼN�U�������6����d�T�լ�;U���TǺ}~���񨱥��a*s��5����\�nu��A=!E��f��ߤ�EB\~�3�>0:@�ǝ~W9���ې&Yk��*�8t��QD�H�b;d��F�����^� �Qߟ]�\
qX	�,��.[�U/� �A(�^���L�7����Dj���[�Ġ(���n��eR,z׍�:0�����2�} [��^fZ� ���5���- ƳdsӲ�z?6��I�%�\���'��n1�E�xK�|<��R�G[���&����ҵ���x:�哢��:�{�P؂WD��0h�"���p@���C��aU�3VRw��s�̶��?f8G2��v��Zp���} ��'SvJ�:7�e\�&�¡n�3������T*���ss�ѹ)�ƄӸ,�A�/�n|���1����R�Jٰk�������a��f�m�G�M����d�'oM������Վ�3�>�6�uwbC���J*ZV\gW�*C�Qt%�f��s�G���IBl ��Q�8~I�7��q�Xܗ ��@�ˣ�XI�tB�G	�5� �C��O�Xn�:|�����.fDx7���p����$~����������~Ϧ?i��cL�p�%�ֱ�=)2�x
\JM
u��I����F�4�P����|Hd�Y���D�`Q������O�D3xP�x�ʭ��ܜ.>�hE�4����AG0�9�ˁMa%9�(��_P�tp��v��Eӛ8�R�D�R�z��*׺j��ٔ�l#$�9����K���:�\{z�?ԙմ&	�M�k�"���'b���Q�NX�꿨�7w7��0U�>O��Fޓ��Z�]p���9B]���Tbj���3,��*��Z���B��mn:>Qu$��<�����E��<�?d�?@��:����i�E�|w�1��X������Q������F�qI���O���zs�ڟZ�ov�٭z�#&Dn�RCm�����AZ�y�n�wA�LD����P�v��iB�Q�8�}��)�S�k6"b�c� 9P�Za!���3�t�e����J��L�tB���|�b�C�
H۹�Q(��W� ��1t�{��桵��׾�d��M�+��6�Z�ד�:Q�Vp	۝�(���c:}�R�*�oǿ��7����E��X�a�{7Ti���My%M���vo�X c��4�ﲨ��tv^����-iy���Ј�L�[�?T�[���u���7Lj�GH6E�^_p�r��K04�b��@�U���4���U�,FA�_ع}L�ޟ��p��S7�l?
���E\���t1��+S�K��٠���|�$oG+�?��7��i���d��� ��Q���_S�d�Q.�+g�b>�R��[��k_�LX���V���۠��X�&��|S�-�9���SS�����B� z����+�pe���y���z�M��3}6xhq,?�Ӱ�3
v*Q9�~��}W4��ӳ�=��H�~�6Z����V�#�y�b����^@�V���l�~�����Z��G`	�6�6�f36��������HW_��ﵗ�1�$�Y���i�/-d�3�����Ilq̑cB�iȁ�Tb4-�������Y��oY��'�sp�3���D� ��z^>uʒ�G���m�%����t<B^�y틗_�/��'�f$�Ⲛ�ͺ�U��eru��o4�3L�,~LO�������Zu��)��~#U]�qZ�E@>�J�D>2�����$�ke�V��#c[A4C*�h���&4`:o�Y%|��%����r#>�Ut����On
�M��n�h�Og��/��Ӭ6����m9~'M��еe�W�3��*2*����C�is��U-@���aT�G7��b�N���o��١^�NX�u_jS3����3�X���Pc��ۡ�b��7�Ɠ1eV.bY�9��h}�07o�o�7�K���9heT�~A�s3?ܭ
n���X6*��r�Y�%�����\�s8�He���f���Sx$��S����	,�^#���}J���M�(҃5G�?z����"���Ǣ;��K�u)
�K\[{��+�r�L���d55�8S�˦Q��Xb�"��۸]����}	�NH ����V :M^�¥HƩ��*�Y�j������M<G_�-����'���Do���İGBZd��|њ��͔�W������~a����3�O��D�5��������<��)c)�a� ���hVc�Eʢ�.�ٝ)�/�'�S/�6IDDR���!���BmJ�����x�)I�_�~슸 ~��C@u���O��W���ޭ��'t�峽/:��aw�4a��s�A�"�,����}K�i3��:>�;;�"W���ʟ��,�{�lo�*9v�����x0Dnl�������RJ�Kh��Y�o�h��.7�V�ૹ�)�ܛv��]�6��w����\s,����*#Ų��tx�F]L��Y(.�����ނ$⚪N]ά�Q�;	%&;�媪T�kb��+4�J��Y���ohH�[�^�*-s�.��U��5m��̜]�n���G�+ߦkZ�����9խ��q� �3�]��2�s�b���zjX����\`���H�a=����K1�l{�E��#C��-4I�␴{�ْZ���i�%��:���6�lW�4N���d��yS�����<"�X���9��x������.ŔO(E����BH� �d�e4���-�u-ׇ9�������:_���G�vTA�x�6{K�u��b���j��H����݀�����%=�����=9�v�֠g�AV[h��(���0ʞHIKs���1�m\d��-DG�*�s*gdEӇ�˚�r����>6x�q��ɮ<"�Q��D��1�/�y��i���>}x���WL�B���P4���,On�dWd����$�U����I�M���N>�
_M�z�U��=�}б/W���J眺�[�x����MdcO³j��rA@���}賩��z���eJ����}+�67nE��ILxIܓ��p�c�=��bjFoQrzO쓣4ku����d���Ly�=�}��,� �c�Z����G��>Ԑq��F`Ϝ�����@�4z��C����ۍ�"P�푧cS���'���F ������WJ(\x�\�%p������JI2�Ҋތg�n��+�J�C�Sja�|�'ɆTI2������PGF@���E�]7�G154)�g�$��	����>�$m=�躹;��	��aȖC�-�%�����~0�T�kN�Y��2��� C%�t �W��"���ڻ�{6j}���C��o��V��a;��H8�l��q�+�b�k���?)�?�X��S�|��#gJ� Ls����bn(t���)�g�t'�<z ��y$ƞ�K�{pa8~�ZH���mJ<̪f��N�Y`^y�!�����X:�����r��Q�ǅ�T���X�P,���7�	}+dXK��niqy��G<3$��{ğP�P?�XH�7G�ɗ3f�~ľE;�������T�ħ7�O��G�2��S��`ѲLL�f���opn���,�.,y;y'9E�G�),x�K�ߥ���)��Fӡ�ޑ�HbH���O.�F|kY�w%N��i�s�G�\u\\o =/"���tlX�������4���l#�0�+~N��WI[J&Ε�'�R���Ј[.z���N�B\8�n�x�6q�	�3�bƊ��T��G�[�msI���χP߲�c���U����1�I�H�qg�M�D<1D��}�Uw�62��ę�!xe��ã�բ�?��K>�z��W����!�j���2��!�	�UI�&έ��2��X� <���AmP��������E�o�[�Jh��WC��
�7܉iM �����Ck�
N�:�ɡ[�<_�KA�К� }�����`��I��!V;����CP m�䐮��/D�B �B8�� o.�ɪ�A��̏�~�^̚��'��.�j#?B�i#��뚸N�M�-l?�
 v����X��@�ԭ��'���_��|�?+D$2�e�|��jz��-R��_��B{S�p{+�*C2��c���G�hi�Hy̆�T��]���@R�ڷ�zI<,x=\�uz�7s����g��Y[�� ��@����N��qcY��
�+%b����YǏ��9���-�J�ϮA*8�U� *��8e�*�s+�}gx�`B*�s��Cy��!\���i�}4M�=-L�����0�?	1k����4�P�=�k�%Љ?�v�:y�=1��4?4�_�� �|�Ru�~*�*u��M\�}Cث��	�]����ۈ9BaS��ٵ����@q�@58=�`Mcꭖ�����{Qf~���;�pPR��Z�9�:[�:в�,�yA� ��9W8��XlT_]�Fj2�S2��&Z������WRɕ�+��z ���n�-�i�R #d�s���QS��8
1ɓ�B�bpgwΚ��#+�z����V`��Yn���s}��(��$!Iv�L�ۄ�Lo�I���� %���j�=^�d��y۠&@��KnCN}ϳ��I��s�p^ �g��38�H��5��1�x�� ��xef�8՝�(�� V� '�[���n׼_�A��՝�d0�Y�*���"5�J	���,�<�l(s!�ȵ�����`y�����b�xU'�Z�S��6w�rc�Q�߹RS*Zi��ZU[���1q`]|��&�}~����Y��iӈ�}kS������X}� v �uC����(�QJw`�!�x�čh��6��Ķ��y3�CE�Y�����4L)g
�t0��Œ@�:�y�x�dn{��Y|��3,���o˴/g}��c�1�q�;�ʦU[٤�ؙn(Ƴ�;�rϚ��0����n�8�PkW��n}�J��֑�R��),��&؁�@g+HV�Ĺ��u�݁)���G|Z ;�3�����|QӪ�a2[������R=�/�㇞c0ҙ�.B�;�k�ASbc�
��Ik�=�c����GI�֣�A/H�SF������f�*$e�����OĠN��f4P�e���3-�"��b<f"<��8^� �o]��b>x����7��F8�>�v�3���f��4\[�n)�~��_�c�*oM����r(6�:'A��f��� �>Hi��)=%�P�Y{�:G|��C����߀J|[m�S�Qj=���\��4<3O���������}KF떋^�Iї�'*6� ��t����F�PtF�c ����ri����Q��t��k���ШO�М�9�j�r�_��w�hF6�X������/�}���mG�*Z�e�DL(���N;�>��~�@�2�]Y�c���g'���& ��mv3J�;Fb-8�R�v&��}�i7W��r$��Y�-�=� ��g^ g������k��">��`�>���I/�{�����ߢ���c`)/���t�v�仢H��vc:O�>N�*Vma7�&��/�z-s'�`��& 2s��S}<���5����>j�F��%aG���� �L&ƹG�rυ|��h�`|����U��ےW��Z� �\�g�h�f`�Y�tp���P)R����r�_h�9K�wgDi�V޾��W)��Xt�Ɲ�m�u�t/}�����(�I��S92w��M㸼��9�NM��ZB�H^9/����L��X���"���W�U\G����{���y|&̈��V��!$e�&��Ȳ�Qh��z�s�Bb�����K�����N�`��<O�p�3��I��#4��C�Fs0u�1#�x�a��
�С���?V�ӂ���+]N|�t�5ʯ='$l��O�d�����n	�Er�߳F����)��/Ĭu�i���\��0���ɍ,-����R��I��@�����aAA��ecSb&�ɣn�f�`�#����ZA��� *�����sݸ)����J�Md�\|υ�B�L�4}	(�[8����&0���x�}�������+�#	E&�����e�to��EyܫlC<Ď�����D��a��0d����*r�����,n:�I��I�FT﷦D ɉN(U5���Wԥ�����ԫ�eҟ��y�0×���n$�d>��㮙=��dK@�kޝ��8��SB�x��mٰ.������W#�fp �-G����ww8��~l/aCf��F¹�*L���������'D"��$$+nFKK�l�R�fI;�0
��g�򃵊�.$o����W^�fڌ��/�U��x	�ݝ�
�b���m��#����k�7�%�v<>;�p�1�G���A�x펌� ���a��t��-��Or2-��:��X��ݢ!��wq����'Ǡr7(�_)����?LZ�ϗInqa�A�	���?o�\�$�F����/7��Ua�S	��ڛ�H�F������Q5F�a>�o@,3�$�nĔ-r�s��#HQM�}�H�C�#5j�������uN G����ab%�ud�<��p�������=?	��g���>�V�@�o�F�1 9���=CM�R��(?�{�����:��V1�g�N����28a-�v��|v"�	by���v���~U�B���b+w�/��=ag�T@!&j��]��S[��ݢP��S��$l�/k��ƽx����EeL7+ǖ��X%[��*���d�������;���r{<�z}A`a_���͞�z(R�y�ݐ���M�����)��f����Z5����[}ɣN�bb�w�qDs���:�7ngv�n��_q�Uu�?/g��П;��uօx�;g-l�d���Cf��'ٖ�i�b�#� �^ď���V��Y�;O�_��g����	W������cbw?N��l4���m���uݧ��[�E�%�/n�k��]��
JšыI���ޅ;����d��*z-V��,�(�E�S6K=��^ɍ� �UN�A�,�ݛ�9��ZUQ�z�90����]]8b�A�����
��c�-�D�K�qpp�%�N��V&I`�2���,׏��v��8O蝉L�1�J0�X�[c�F� �W��U�q�<�HĨ�c7;�Y�
�T�Dk_�]`���bX*��[mԶ�Ε�S6�efwXh�,>J��'}�ln	M<Dtn��$c i�h��x��ő ��*���ȋ����5m���4�Dg���D�`��u������
 �诚+�Ն�9��~cl�	NŸ�-��tp.�#&���8A���"��#��s1'������L�E�[_����*��(�h��=�$zN��S��ٺ���(\���t��<��s(�^o�O�J�Ѳ3�Ƿ۶Z��[��c�t��_�V����,�y��oϋ"���vƓ�@-��� ��S��26��j[�p{��cyF�b��(���]��(�^�� {�����<	V8�Ƚ�60��;���Th����N�����$Ǵ7�f������D�'��n�'ۄ���M�!�!>��*�C�59��x��SE�l��Xt?�(�ǯ����8�~���齍�g�k�c������*��I�2��F�/. �����h�7T�K1�w7;�g;��}��8�op�g�W���6#�bX���I��X��h���p���O��'�Q�{7(N�:�[� ~2ԏ=�OF�l2��1�I�0� d���^��05_������T���.�5�������i��B!l�t;��}�ͫம0Ԉ�0b����[���ʁ[mKa�DݫS��t�e����'����)�sd��sL$γ^�h䐮�e�+���#{��6hT{��[�pb�>����o�,��k;~0�K3qʇ��!�d!��N�F�nG�f?R/��naN�,���hf'���IV�eȳ�$X�aYw�S0�}��Qp�����ѡ�}M���b�h�n�k����s�J:�c����06�2	!�~.����$&��t���#O���'�'��q�<�w�"�l�p�!�1K{�_x����N!�����W�F!@hO���p�����)F��18��s`,z:^l��t����P+m�
�v���Ԛ�D$��)���":�O��X/W	j7����U�A�� �TNq���Y�W���&���0C-��x�k�O�t�&�m���q>Y!T(���c��9w	����Lx�=g�Q��.RN���3��Sz�d��h~�u��x��<���I������i���.��}�ɀ����
i�g��.�R�GQ�7�-+�h;ݙ�hN���ӎn�Ų#����#cK�&\_�~ֺ�.�;�Ap��Q�5;�y���䏹�m���|�q��g^kH�<���G�$��9���'WG7!��7�:'u�6��coxo�����X	�$&)W��[�I��BI�BO�_(�G��qA��V�ī��y>�ţ����z�=l�+����	�Ť� �}�*��+U-�qʭ�:8bq2��'��� �YE�|%�o�ne�T���/�,��ҧ쩀s`ГiΏ�Y��*���lY�<��ȕ�R�7�h������ ؜WX�,>a�f�&���Sg��hT1�����v���i�FV������V���煥��0�Z{�gܸ��ò�g��
�%K�(�����)H�i��`��q�$�"��8,g1���*%��M���NcY��g�]dx�%Z�
��Ʃ  ����n�@�mv���0��!�D����d_�(4M��1����W	�W/?��[Fw�*�.LT(��)�!�1��<ނXx�dPv�Ϧ8	�����.�m�����(^��C��7�PW[���%X2Z��S)�
�P9צ�1'Y$Tt�ш���;W�o'�K�cGo��h��n�d)-矮F^�mB�Ex�"�zc��0p��>1�gR� p�$�9�W�'G`�$��HoТ��!O��^��w�����2��r�x��-:��lp�0�YJ#��d	:���]F���� �8�9dg��?؛���1�#l��]�7=bͶApEQи&H��܂��H�N�۴EM?7b��98�Ùƣ߂� 7�s�E��;�Aؾg��Ή�co7�r����>���+��Q�x������D�00���W�]GP~�����()L}ni̺ZU�ҧ�Վ�Ѽ)��Vb�2��}ެ�78vH�g̤���G|�O�ɵ
������r|��Jv��%��j ?����&��,��x2��/Ï#8�XJ� ѯ���O��Wu1÷N%2�����S<P�J�ڜ.&�j�2�.8_���.6!����'��-y�x<v�^�p�aKTI+�N��=�T��B�֣��$��Ÿ�y�چ+=e؂Z���G��b�WU_d&yQ�E�I����� L��A^O� t!j�?�{z���5+�΢�h�v7�����9�vd���M�/Tv�LLٚc>zO}댌���=�)�'C��*;s
f���ݴ[M��d1�yA�3�ʎ=RpG�k_��U�&�m����j��C�!��zE[N��z]���Nv�.��;Y�Y�R�$v[us)�!�Z���R��W�P	$w<�#�sU�h�KjJ��7�gZ%�0�2�{�A�a��da\~ӿ(b�s��F�%5�\�5zW�������p=���X\��CBfE���$�ŷ�il	Y5l�0k�ѯ�b�y�lT�O1g\`ޅ2�{�����n�E��]��xR��U-��;��:mjdTK�p�/Wh�yu���l��b�!��&�u���u5�oo�9l��R���kv��_$� ��>L�s�֓��T�P�OW»�32�����{�&򌧣�,���K~lw$����v��4ob�e󦰘��::c�W����(#ˈ��ą�J��N�\�p�K�1�M��k���ED���W��-�3�l��u:̍�{q?b�`^����]�h�K�v�����!�jB+�[�r�I��Q�u��z#rһϮGH̖]�O�*�%at|�\���|]�g�q�$�������M�INzal�T0��}��d'�åyiDt�V�իO����_=-�Iz�KbU�$�vB��b�	�<��!%H���5���f�a�
���JsQKx��[ݹ����=i��тZ
q�����FJ
L�_N��%ws�ɻ�Q�_VM������5��h����E�a���P�`�`�Hy0֛)�Ƶ��[�F\
"qw�m�&�!���2�h$F������E�H]�r�S��o��V�$�M���J�9�:s�Ǝ��d����2�������;ϕ_��~��`�x^�46b��>^ ��R���@�Ab��?9's�����
��D7 ք��Xƀ��������BQ�S��N[�G,�Ϻ�+�G1�0�j���6��/��_�?�]���p.�~A�疡	 r���v�.�}�4��������.�٧��mU�c����@�#xh*��ЩEr���h8�t�y�-�hnd�{g����0���3��U�y�&���=�	,�Zw��R�*�ٿ�>
~+v)Y<��I2�� )�q&�kB�^���p����R�~ 8�3i�L�ս-���B{v����Ư�F���=��iQRh(��r��28�^8�o��o_�����Y�9w��u�YG�����ƿ��a|����B�Zl���X��)�ts�8�x�,�W������Q�M���X�`�㱷n�\����^L-@]�V�F�+�f���[�)�B�]ȫ�������p������LyDU����2�\��[-N�>������jl��U�#��}����Eڣu�=CK#E�C�*?�����5�8��B�$K5W�!M))#�8��b�x$�����C��5���X&�k�:�p�� ����g@߯���m;e{*��Grt��odū�9���e7�z�J�X "��z`s��tx�cf���{,m�-Uo:��[�t�����������x��֥~�bқ�r�~G�뚲,�����f���$Lz��j��&;X��i�	ӓ���$�i%sY�d��{tc�`�Q��H'��@qH	j"�B�t�	�z�h�+�Q����g��'���r�F�BK�u~�i� Ŷ���bu5	h П!F�Cj���l��q���1fa�B�;Lc�3;�Y���.�=��lÇoa����Iq�\y����2
�-�S�H/x���W����n�E���>%��b�v4�@�I����I���Ũ����O��~#�4�=��b�c������^�OlZu�μ�]w�m�g:"|VLg��ou\U��j��#3^ISr��ԝ�gNA�`���bo�O�Ѝ�
�`���G�2���)��R�J�8W[m	4l��.�%�N��q�D��H�6�<���;��<�f�{O�'����W׫ý>��u����K�G;�xRa���s�%�￳� ��Έ�{�
R �*l��w��x>���W�I=E��XI$�ON��:O8T~K��!|�F��έ��=�j�|wbc�z����$�J��-��t|D0@���"7��8	�z�u�)}�%�h�{=b�'����:,A3\,�bY��Smp�甛�Ӽ��,�rsGh���ђZ�ڟ�{���-�'x>(s�EZFA\�����-*�VJ�c	}�v���g�ׯ���o9�o��~�/���5���u?{�=���O���+ˡN�M�*��9,Asu����Pxcv�F�QhRp6Il�l�Uvr2���:De�5�q絗]�5��"`�#i��{H+
�S+�5���yA]�6�p.�]f�m!!!�_�d<w�P�`�Q��/�|G�6�i��2�)�ޛ�ͩ���1���.`b�/���W�y˾�]�>�GQ]3+��c�3E��ݱ�Ng�j�T��l�0^)���u�j&�ҵ���G����1�^&���郘k����Y��!����S�UI5B�ZAB@��e�\�dc��ܧ|�����z��8����Qh�*~_��Ɠ�G��VfaG{�
B�be�F�[-z�PcBrҊY�dE>/�~k�����#�U�>,��@�V7h'�ܚ6k�S�^dhWǕ��Ϗr��>���s6V>	k����c�a�i��h�T�l���8�(�c��%���9�bxn��}3)$��g�c;*�pi���n�[O���=���B�+G�鈸�e`;�2d���-�=�hn���߈�9����v�|� �ؙujY� hnZ���*�*���R����I̓����w�|��6��N��O.�ˉ���7���n�ߪwk���B���8�`�c��^�͍�,S\�-�|Ë�-*�_�0.�9O-}�lG2��"-�O!_�w@M�����6%-�Llb{�B����Qᕹ�2���uD����71M`4%�^P��z"b�qf��ŶtU"	Ĳň�R���6г�lM����2�Mų��R ^Џ9�45�>�AQ������P�5ѯ-�� W�Rs��ϦNf�د�L6��94'��]� �6�K<�L�,��/���0y"J)��o-F�&��N�=�2"Lܑ�T-��-'{�C�p�ǔ�rx/�"&��������>ɮm����YN��}���GVx�*Y]��1��T��X��_o>zC�|ZW���-�.����S�����.�	�מ[�Z�����h`�<"x�	���C_0-��o�J����s�I��XO>�ft�_t�Q�]�L�#,l8��JխC�����/3\x8A���kޡuK&�� ����w�r��v:tE&H�<9:�v-�\%2�yI��W0�,�(�:Vgȵ�/��T�2�#dU��s	���7fU��LZ~�?ש1jN)EG�$U>x�=l-���=m�������1�L����t������0vRdW��2�U��J���|�hFc��|L���!��&~�
�m���h�r��%�����~������N��������K^F-��za5&b����Ӎ�= ���Z�-�vn����7�A
k7|&��/��������Ɨq^�|tX���l������d�6X��3��8��L��7�H���%dS��Ǝ���V��}��?L�������Na��g*Ba�K#;\���v's��D	�X�����X�c�|9x���TȰn���Z���);�b}������B%T�z絕�5A�-�`�N*C�����k:��A%�*�fP,0P���(+�ͳ�w�C	� ̤�m���s�<��<��b[vXګ�//�U�	�6�4�G�iG��Y�BZ������Q��j��?�I0Z�i�&���D�̷bd(��sH�~@jaaq,�w�m����pE�1��X����O���^�>���-�yӈ|����jLQ�Y��Z�)%���5@�.�	���*��T�:h�����A
�-H�? ��?����_�|I��ͷ���%�I�D���/�/�����5�th��.�����=�EĀ\��6/r�%#T�����i�P2E�A/�������^.�`��I:�O�^;�:/;x�����X��+	"X��B��8o��SAёx�[R��%��G.�w�"�o�o�8��k �X�J�ѥۄ�,��|��
	������c��]��+~�������&tL���v�4�Q�Ӷ�U5D�cQ�V�v���2�C�d]%F�o�n
wN9W�ު��7�y70m�C0�Ie���^	��>#p�_6j���-k��r���R��o��.��zk���av��Q��"p}�2;�	��E2aS�����ҿ�HL�.\}�DE#�zG&��hJ%����@lr�]5�Ti�3��.�N.�S28�~��?&��������|!��Y��d ����TZ�5<6�-Z�4�N�koAEK�(����E[�uʬW�PG�F���h̿'���mp���\�i�St�p��S(n�dB�d�G>|��Ym�$�@e�K���d�.��LVS��s�u	9�C�~��ޘ{�٣�ה�&�Ǎ(�WTP��Xߒ2�,U��	�{��^/��a&�`|ff��ݮe�0�F=\B�pR"��Kr	��S��~5{�b�޹�X�Ъ���_@T�q��V��\!�9���(<���S��	��ߤK�u�%ٰEI�j�5�����{�Q�u���4��P?��U�G蒈Qc�ul�:��������a��\N�T�hC<�@cc��� �Fi1��|-����Q �T(~Ɇ.���~k|��c��h�]��=�5N�qc���H]�*�W>�G}�h��ô��Ƹ񽮫���\3n��o��Ձ"�=�54�%�O �HA� ��e�=�m�����B�U��ʏ�r.� }k�Ҭ;�w9aB������,���>sdȘ�V�M^���ҹH����a�1��j��@������s��o�ϣ��wLZ6h׮�S
@-�c�"w��qO%�&�6ÔY��M)węԖYw1��t<�@i�T���ik�Я2̻���>�;�?:�t�Ŝ;��#�g2�ߤF�����d��I���i�Y�O�g{��s��fX�?�,9��+d�!�TG��Q�Q`��4����7��?�M`����Rp����T\lYF?-21r5����Ok���ں9���!4O��N��c=FAuF��ؚ�6���
4�q�
�K�0��{�ұΚ�A�ϠH�4�)lk��YGYu�x���v���z��G�k]v����{q|��r�7��WPN���"�e���^����)�M?-a��"���{]f"���H/�H�c���Z;L�$"֦�Q��9�������}����c`�9^���	��=Ĵ� ����/sˋ�&XV_s�g{�:,.$��Jz���T�q���I�cփ��!Fv��p�Q{�=Sְ۵<8���3D�ei��$9�����<���`}$�ȗ���(|T��r������as�8=`ay�S���G���(z�7Q;I<Fn��M[��,�n�g���t���JM��A�|�$�Z�2>��eˎFtC6�+����Bi���ܣ1|�
#)B��jq&Z_�3�=����~V1�o��;�O�jʁ�އ`�4�UN>���YFKy���.-9`�ss��_�0�8�ol;!JƤH�g��:U�4V�D��Mw�����<��(_�S]�O�)�m�m��sR#d�A�Ih�"������p}5�r��Ȝ�*�����2~w-�c3Ģ�B�"��8<B��ۆ�I��8wF89,A|���ь��Y��]��6Wf\�o&+���&�Ggӈ_�\rY�M��'�4���*�E��
㸡푱\y����%�Ʒ�C���սe�%&($ ������VT����$��_�����>0R�JAv,�8ҡ�����rb��[���y���èW�K���&ذS�Fy��,�m���n5'�O����Eu� ��;"�	7[$�����uh����/�؍y�BQZ�8j�2f��7YЛgaC�s^8LW���Q���4$��nFd��f�H�����^q>c��K7��t��0Z��Q��( Y�`N���٘�@��;y�BV]�=*�a�x�Z9Z�2cdZ��������^�u| 8�D#b]YZ��%��p=BK�
��C.{L�b�4��e�CL��/���'7��M����������[����+�!.V;r�FB	F�����e��ŧ����#��ͅ�F�sx7'vV����	�pǆiN��<X�nNL����nU�1��;��+say�:YPQW����V(^5�$jȲj��CN���ޏZV8��`��^���Y!�a�U;ģb~EE�R�I������DQ� Rh���t�s� ԯKZT�HI3��;�(��&Lm�}V?[��[�*G	I��t��*���M=���^���۵<���lWT(/���J�����/����%�WN�2����j���K<���H~={"�X���w�o�Ƥ8���.r����6���=Id!]��mh[��SU�&��F)��3i#��|������k
���F�6�
z��As��A"��c[���V�=@%"<�K��ׅ��F*���x��vF$�m���	z��L��}E��`��g4��;:�j��B�5���"J���vLI�pWU�$5H���Ct�r�Ͽ0���t�N2�O1����"os�R�^�ړ�
����U"�7p8Wnl;J��/;m���o�H]�ZP����)�bxJ4o:wm�EǗ��f)��o���z�%��|�qo��Ta��;[���*N�B���d\M�z&�Q��ȳ��ı��`�WA���e+�͍����o�6�<f�[!��`1�Yc�D��` �
:{����]U��5&�OY`���B��4��)����hVc��i�ݤ�X��,=���n�)8��_љՕ"�N� �K��aBj�j����;T�ѷ�҅�!���gx��`mHN�Ϻ.h��&�zt^@_���1��ALù�H+����w���?����S�+��G��[a%<�,c��h<�/0h^TT����"���/g}�d�¯���Jj|�����c�f�����>�<���([��L�6�KlN9����*t���$�~&�����M��yJ���%�G�rgO�^UX�^���A�{Sh���`FD�U��{+���M�t�ا�������L��2�!���{匷��0�ڎf_�4�3�꺾 m�fE.-[ШӅ��z4iVK�>ڢx%}/)�	Zwh�8x1ma�%sX�I�)+��u��\"8\�xk���0,d:���A�Oͣ�����x���T�?����J�4X/	>(�䉅nc�)
�+����N8�'�%�p��gzX"�������#N[�Zo4ӑ˙S�)@���/~�ZS�7��
C)
ǎ��������E����,˓4�� ~zo�,#�ȓ�-�`���F�X�K�&<��	�5־�xkTz8���*� 
B���3�՝�����8f��1�M�>l��+K��� �\�MQ�l�Ƚ*���IG����{I��r�(^���(w����*GF��C����������� ɤt1_�n�fݽ��إ�ګ�����>�}�5��Q�����B	^��fU�Y�nD)r���=��K���u�,�ŧ���[Mʰ�\�\��l~���W:M0�OE�����zS����S�e�;:C^鍟I���p�.�37�;����'�b��,%.]۹��E�+E��C��mY�A��]r�L�2�,�6���I,F���=����`�6u{�y����wr$���o�L��C���8�^_Q�fl�BH	!_�}�ߴ]0\?e�{����p����H�|����z�5��K��T˿bh��חj+�!���m���%7�XC�$�YW�����AI������6B%�	j���-E�V�_�Y~
I�w��T&=͙Rs�����h���O\�S���=��qNY23|C��]��s3�`�$��N1#�!�C�=7�����_1��\�Ǉ�\�`��Y��5�p����R��������+�<߁k%#�*goA��M��Xx��C�%��l7A"܀m�����԰M�p�n�ip����;PvY'�*�&�W�Q�Rg*L����0��u=�\VL=�0e�1�W��<������R�
�s7k�?��TN�>�aa5j��	�p�i5�y�A���Q%؛�	-#)�v�R��/>�;:ݮj�j�����a]a�+r��6 ���e�V���(����[�=�f�ʦh*��%���!С�(��-YT \�,�C���u���[�L���m����b|�/��(EE4�W��(�l��D����g{��^�e����쐌��L)���f�tS������N�XdPZ�c �+��-%��j��Mà�*!�a\h1�*����5��|�(�Z ю��P�鸨�-2B=��.��;s�!��W�H�ɠvr�"�0�Ƕ�ڵ"��C�u%��ȕt�m��;���'�^;/�y�K�i�l��*��|��+O󞆹�˶�jؠJQ����Z�Đ� 	��9	X%�sV+`��=I|߇qI���vF�'V��To�������o��B��2�ËL�bA����@��U}���� Ŷ�9�����JN�$�<H`��7��� ���G�!{���(g��5�8�������>�g�H�7��SYn,e��y��	�i��%��p���� .���j=�����OV�r4�EՆ.��;d����U�����e�k�..��Ay��[����%�<B��&�Ⱳm�O
~R�@L�x���K_t�q���{y�c���C�j�S����ˑ.����)�/vM��`�UՂ�N�<��ryKG:��J��}\�tP-�/�	c�x��7H8�'j�^�����`T"t����Sx�%�,����J�.�⪝��N��:e����}uO��U:D2� �FG/�D2�:�J5��Z����4��u/�8l����I����`֢��ĭ�;\����Q3�vB�E��ӡ�~8^x�ٸs-���r�;����}�����g3�W�jO��}��M�D)e
e�N��t���ؔ��L-l�����h������}ۂ�4��%�>��ն
�pd.@������x� ϯ�͒�&+K��B�+M����l+�,!��瘽�5(`�9��<��1'�〞$���ͥ�P~���z
O�����vo�5���O��iN�	���wyZ�S� ��f��i�Ԃm�/�<Ǔ��p�E[a�$����T(��I-	ǥ�| ��(!.G��pr~�އG�c���o�ɋ���#���*٠�r��۰p�������`�¼���0��abBYUd�e慖����d0:�)����`{���3��ե6�is�o�>���Q�٩�#Y�Mfik���=J}�Q@j�N���A�^���рԳ�k2!����Yb.@F ���a膔��������̉���Μ��S@�q۫��y�l�I��W#����E"d]�i:��|��c�9yP7V`,2����L�ٙ���@�GO�˾�Nx��'�M�4�����faت���$Y���Ӻ��g/l����KU�C�D�!{�>�@�`���,��9?E��F���HeGm0�A�h��w���B9*X2G4��n�g��`1��xQ QBj@q|�U���&���[��Z �?h}Y���T��/g
H"�B5� @D5�qTDf6���T�\���Ƹ�1>�F<�=BpJe���m��MvH�_ampz�	۱f�.Y°i��m�*�]���>N�����y"zX\�ɐҶ�'�� ƕ�"�C��0���=�y�;W�ܾ�y_��l����z���m
����V�5Z��nVA��m�	�4�:\#�o%/yxT��]��L] ʩ�b�>�h8�%xk���m����  �{e�~�߮��0;���r�Mn��%Q��,�x�͍��=��%}�6�x�+�����eaȞq�^��V��n��暻PY��{$\�pV��3��/�6 �B6G�1%-1����z�J��Q�}^|sx�rn�O���<6����;��p���}��f�q����A�sh�~�rhsf3���+�.IPL��r�p%��`�-��Ӽ�R���"ֶ�B�������ox�b�;���"G3�y�R_މI���b�B6�y�s��<��t�J!d�-n��U[}�cb&���#U��:�`w(8ְ^t���X=���2����j���{8��_�y�I*�a�������*
�(�
|�t�xt͔!*Hu�ά�e�\5����y�x��[�*��`����w�e��(�=���F_�v(��&D'L�.�V�J��T5�=7(;��F���>n������}yg�j��0�&��!�
L�(���dD'�e"�G����w�SvBc7��H� ���0��) �&g��I�Q\*ZA��5�*����z&�:q�1B���wr�������_�N6�G�b�`�~�G�����x��*z�z�z��,9�8m|�Y�����NO���E^JPRa�4��~e�� /����H˫��:�s���q����k��l@@�	!}�6���V�2�w�L�E�}#o��ZP�TC"�E}"�*��YK�� ͡Nj�F$�`���j=gOOG��p=�R�j^�Ϸ>=�b�0ՊҘ���2?|AC`�>r<��TY��C9����Ȋ{��ZK�H��3F�ZXj:轅���>\M������}�{m9���@G�|�6^O!;\�;����Ύ)�ǥ��*>V�?���J]�:�0�g��g�,@����H2�Iv��K*�7�Ҫl2r,���|#:d@_C��p`^k�onS��S�N��]�l�͘��f
�S}���Exg���@bFs5Z��ŗ47��v��;-�����S��mW@����z�|�R΋����͒��j���L�YHI�.��P�R̆v��L-�V�8d��Gk��Kd��TaG���� ��Ⱥ]���YQ�f�g���3PϨ�i��_G��Gn��//���ѓc;�V�^�;��D�{^�{H���"ߎ�I���5h��7��lKF��[�}����K^� Pi.f�	ͪ$� ��/@�^Գ@���o��1�	��j7�-#��.�ys��%����S?��4Pa.c^i�߭��n�ړ�<9=��5���!�8���؏�"cY�v�>�)�m?��X�P�Ĵ��QN�4+B��rÃay�A�M���e�}s;��̯��!����;7�++մ9�s��ph�����w7 ��@�P�� ��#v
#�I?#T�V���ׇ�[����̓���a�7�@S�C/r�C��{���x�t�*��b�l�모�n�%=p��x�`��n� ���ݶ���4��IE��?�r�x�:4���1�tFA�~�	yER*-Ka��.T`S'��l�q��.kJї��'�q���ֱA)W�<����y5�6թS��J�1�zӓ��¸[������\��[��gZ�)�I�V��1Ғ�5�t���j�!sbC֣P∨希��W+�8�����|Kh�6,v�?UFĻ��\hǬ���*� k:�M�f��71�Z�,`��~��3����7W<է��;�!��,�э�U��4Y��Y��\z�cB���uJ�,츥��a��Aq��7�%��D����e�:%�jzl0/߿�ᦑ�*�]��#ZM�g�7���}��r�>����q�7�_q#{Qƒ�r��������fKq���/�i��`�r��3I�$S�Ʃ���1��XB�ǊQ�m~,��@�ɱ��S30�{�O���O�/���+���Kdø_)D;�}0��S�+�9*!��B��%�
��xvB���f��Z�7�z�RO����u�p��C|�8?���e;�I_3Ў ny��ݶ<�{�"�;��dX�T��YI�nFeY��y�e'���Ro*;DހN�яU�>�5� ��G���#�WbC�v����1+'&�;tr��z8J�?b��Meμ�5��"��w>�p��ߢ�|HM����'�>,�����s��>�l��n�6�q�}\R3e��Qh �c*�_bD����̀q�*EUp��.�'��y~�\�,��eӒ>��9?J�G���IL(� ��g�u~^d�J��*ŧ彊\�$�-���͇R�s�ӵ|�ӝ���������{�����g��>�k�J�QޥW��O�S�iq=��-���� }p׏\J�L;2�b��9���x��H�,(�荛,�>{�<�6��*�,%�aaP�K#�3WC�/��LG����^�����a��j�e5��3ͯ�'�s9�a�L�K�[�����@�n��)=ϟ��є?�� �d��U��D�չF`َId��b� ��B>7Ɗ�œ<F.��O�'�(<j=o3H��ʐ�Y`l1�1x~����Y���/����[~=��[�1{ˍ���Ĩo)���bA�<�(� vr�99��-a��#��fQ�ҁ��6VmI7�c�nb*�����B#�VPZ3���y���zZ��u9�'�<��ƍ �g���2]��kS�[[�8���IZ� �X_���Nt=ź��(�Mx�aa�C̯'�z�cK#����j(S]��`��x:9�'�������#O��0g�L ��x�R�Qi(���@���UI�O�����'�u���u���{�ܤ���X�V�}�!G��3���Pϳ���)#hId7��q��J�qX��\Z�ܡ��"06�Ѥ1Ww_SAC|zG����ml��*�?p�zk>�F#�̥(��6�1�I!�P�}�,c�Sv��w�j�E��˃���<VG��#:xZ�.�!�2����
o��� ��ϵ�N:=:�%��!'��}y�id/ˎ��~�4845�7���䈖�����i��{mW�|t����%�q��];�t���a�8C���Xn?���_w��
��MҬ��ڢ���{�X0�ʤY)�6�.�k�5���&��":gYڏ21F�b��T� �	~~��b�l����\�v!/Xv�+���o"ٙ	�u,&�w���A�N��&PK��Di/ I�̇�.@���q�H��dGzsYL�����(?2��9��	姅W�@y�{�'c}P ���2�)��Gu����	&�A�ۘk2yUIG��;�\{��x��r���Y4��P���ِq=\͘�\o�x	Į��/�Ɩ�2>; l�U���p#�$|�-�����s�=�ҧQ��J# �_��ct=ape�y��Q=��!�?�2CB���|��#"\OT�?�α��!�SG!,��h|��/l�P�A��F��o}����:�G�1HEn��n�u�l��MAF4�P�h�c�8�����U���?|��4�~���u��o7K��7�t�V/�)!��������R�\"����]�h�[�4�?�w�*TOY�t-�{2����`�4�y�X%����U$� ��PP(�0��Uh�̹F�����^��;��Y�ΝQrG׼�W� t��EN;0A�5?���h�*x`��� ��Wgڟs�.sJ]�7�t������-�*Ҕ�J���4�� F��@Y���Su��(�y"����p9V��C䵔{V�����LA.yH���������^���S���Ve{3��{g9�y��q��T�L�%ՙk�b��2;*q#!ﱡ�:�\����WD��3ȼy����E?����Qm��lY��Վ7,�1u���㴿q�'��Ko�6X����B�0T��=�Z���C݌SM6�k�׃�'�N��E��dMw�I|�������/��!�]#�ĺ��:ւ̾�7~@�+���=��ɓ��=]�np:��ϯڏI������	6�P!M�J'��)�����(Ͱ��Y	�!� I��a0�Jn�/W��mK'��/CQ������a��(���Xv�Pl8�M?ޗ�`4X^�)��"��F�16�l��'�~���Zڴ�L��ɍ3Կ����	��ƈ�vHDx�s��p��Xl�=������LL�s1��]�w��F�fY$bl�;�S�J=��g,�6�ȵd��5�R;fúhٴ+��_QJb�=Hh�o�����6�E��Rs�&��\�w����QD����
9�{US_a�I�����[���ڂ�q?;�I�-|�T��LVc�KS>0z��N=v,��	ۉ������hq�I�%��}^a���Hb���+z��_N�H/���^�����a
w)����M��i�&el��xX�g���&����E>��(�<��Z�K'��?��B���5;�DB�� ��~�t��A���y��l�����9Q�Ld�S����I��fM��4�ЁW�C5�L����KU@A����Ȋ����}�Ϳ�/�4{ך�7fL��[H4�P��)Z >V�����ޜ4U�����f%ɨ��O�[}$f��з��GlQ��ϩ:0��� ��+�j�--<��ƲR��u���R�2���~�|%��3h��,Pxv�6>Ve
7�vam�W�\�#6�W�g�3��ޗG�)FI2����y{Fj.��7������j�O��Bӷ�bc<:(���JID+H�=)�֮
m��z
2�ʖI��j-G:SS�B�"�I7���b��AJ�R�D�R�Q�
������$:�F:i���^u��1�܆%�
����	g�'��u�˪nV?�q���/K������4t�_��1��&°��KIc�pJb��#<{t�<��n"g+�ӷv�$X��2�_�ܚ������P��e%c�O2���|k� t�X~X�Y�CU��
繨\,#
w¾�'�;B{9�����']n3�9b�Z�c��N�ϷFu	��dM�@g�.��{v%�D��p��? �A HZՄ$?=҂ru�v�.��R�4-y�-��:��5�ಯ�G[��!h�X�f(�a�~6����xjW/�����C�S���w@`���y�c@��ZgE7�	끯:�[�.=g�9����,���i��F���=C ��^^s�����$B�(Cpc	9�zafI�a�ӏR��īk�~8���{v��*����F�x��w>!�ښ�۶\�ȶ�X{��py�� $f����vS�-�Wt���!�ꜶDifP���|-+mS�r�u`��=\���C�K�$���h�'X�>��=�F��ƍ�C/���׳���}K�^�E���mO�W��ǋ���ō�`�������R�� r��Lp���� �Y����@�) ��1>������뵶w�y��xH�0�d����2�v�7[�=�D����aJ��w�+4nn��!�!x�.�t�n���d�1zmj�$)<�[)��7K��W��ʌ}�&���oCLS�55!����b�r�I4d�R�q}�	����M��YȂ����[Sܧ#F�6%�7k�}������TMA��/j����QfZZ	�b��3�5�0��i��}��<��T��>rv����p� ���do���(���m�(:��&,#���u�Sx�V�4�ڈTi�}V�x�Ǿ,�VS4�����P���M��6i�� ����B�ƛ�6{�^|+h�4�3O�ry#���"p�'����oۗ,0jt8$�>�*WB8L�V�"��\����������������)����>�ʜO�l<�H땬qwt�\Y$�A�l1�@ʓ�':�;�����7]����>Y�\����hk��z�j|.��7��jb��D���d�^���*7��'��kS��n��N�&�i�B�ABH,X�
�2�Gs���\mt���Z31:� C��뒺nsF�A`�V {�:�xƦ�	�0@���-���T^
����[�#���x��,w�(V�d��ë�s��9�_$.D|ʼ�����w�Zq��G��,t��< W�=*�xd	�^�F������>��"t@B:��d���9��M��Ԅ
�,v�7�����%�}lXK��>�򏕋���G�g����tܛ���L'�0Aם��:;$�B�߭y����/�p�[�n��֬	���S{�7�-�k	������C�6L�盆[��AC�9�0� 5����j�\��ks��5Lp�Lx�����D���vY�JG���Ӿ��B�g�M#A8?(��`u^6/�dh�Z(;�+�qМ��Z��\a˪uN�u�4DǛ
��M�ML����6� �l�S�:9?�t���0Ƈs\+T�a���(V�I+�� �cA_���f̵
S9�u����1��R��ƭ᝺��/ �����g�(K_d���K;��+�L`m�*TD�'Eg�7Ƒ�W����{I�Q��J�3�6%��vʳ�(��N��n®H��C�w��<���H�7@�G���~�a�$P�g{�5 nv7�%��y��B	Z�_XI��������T*t�H0o�V��y�Q/E+��r�N�k#�]�s�v�.꜡'�z�>@xJ@�s��4��Q�	��|�z�]Tt��_��GP�/��ޞi�GV֍�𷳒��';�կ�-_�t좔�P��A �/.����p�gT��m5q*���p��2���y"6�w�;/~�y�E�X�۰~��ߜ*�q���ayx�y����pD?�x+d���'��r	��!3��ҨwE�ӈ� �Ԏ��X.�N�;���d�$KmUL��r���� ��p��vB6�0 ��{����q��N ���F�|Z`�I���l��0j� `;[�s���"�
��v#��0q<KC�L_.�|�8���NV��ՙih�	Q�@� @��OH���Y=���Ua+�/�L#b5��������n�a�(��E��� Ѩ��g��̫�7����	������-����/�>�7�f-	2�CC-b������$���n�V5�q�����׷:VoETn=&���v�!g�#�T[f����������k����q�w�4�$�K�|�^�Iֲ�>^�L0-f_h���3>N���{0C�����<c�p��,n�n�a�\�;������E
w���s�H-�b/�qf<0T΀v�-'��Ҏ�1t¶����p0��t}q|tv<��Z�eC���~ m��ʁ����l�f��'�hE&mG�Si�a^:�x�	.�*��"���J@v}����c�-˷{��Z�^u��*��U�0�!@�x$tVD�-EĹS:�����˂>���S&L;�G��;1M"�����.����~��;��c`�.̥�P����� �;)b2,���s��v��c~��9�r�|.�ogQ�Z����@]���F�7��bC�t��~�=~H&�*���x҃.B�5��e��e��
8�g$�]_��� �}J�2�������!��R��_ͭR�G�k�֛TZJ7��O$ڜ��$Bi��p#Mr�'8�Ԅ%1߱|����g�@�mH�����`=��x����*IfZH���cS.j�m>INT|�(w N4��
8���H�����Y��'Ĉ�e޹e-��ES�'f\�G�{��#��h|oAdJ����	�&Xn�@��Xdj]�s��M$�J�Ψ"0^�;�݊3݅��Q!S�c�;�λ*��Y�����Q̌������n���8zk�;2d�t���x��B�^�_�+`�$��'ISA��)�����^I��g����9�q:WD��[�D�{e$aE��n
�d-�<��<���d�U���8U��[Rck�@qS:���D�Կ|���qH}�
j	}������u=^]\_|��,�LPJ����6YЪ!�2i�%Dc����y���O��ug�*}R��C�>��'jϯ2kk���f?�I�uf��b�a��3%�,�ZRvܗiŨ�#��z�_�iz%�r_
�Z{��eur�R�ə���Xio8� ��jQK��XBŇZ{�=r��q=�7�l��Z�&����YN��H�a��w:��@��`�*�wק����\`e�H�E�3���F�D������}z5f����{U�W��+Esgd�s�?R6ۓ�:MN�\�V�݄.D.,g���'�o޸��7�@ʅnIb�m�������Ƈ�m��S�54� 5A
�VG�-�}���Ej�V����2t!�)j	�����x��9~J.|�i��X68�(�9�wH�ە�t7�|2���X��^�$��*E�;l���(���3>�et*n�-��窤�����s�w�� �_�`}W<(�v`kf�����زs͸ᮍ�g1c���Wxh���i�(�CRT�������0�	u�Ra��%�E\nLK�� �1�k�>�#s�m�/�j5ߎN��6���{�ZJZ/�T0>R�qBJ�ks-ٸ��ҟ��[��l�5�|�` ��)eC̅�	.�~�����P�9���{�񷀚���-W� �Q�v�F:����{/���/J�����}�صi�R�i�r�'H���_��W���M^���D�U_�yq��A�+���SB��O4���m���5f�C��.iB�'�1t'��j�O�=/��\�v�F�V�=x�}�7�
j����G�/�_�2��H�Y�(F���?��lW�K�~%��#�H=�t0"������3~�6�g��I�X���C� $a��?8�V���h!��2�����;|C���L��O/��GK&���:��Cq��3���cZ]̂u��<T[&ބ18d�jqǢ,J�9QSl��qk���s��\&����pw#��+WTla��kiI��Ø�N8����<���5���u���Z�r�(����<��Tw����؀x��c�2m��%�/�E��"�������j���,�)�6�A����6.ݝ�mܛ�ŁsY� �L�RU־rڜ6p���-(|+��J�Qs)�"$����M��Q-%����ί��,~Eܲ���B�_�oL9�ȷ�d��,,� �(�mcI��={帏ET.)x��č��J.�!
rYS �8�
X(W�[���t[	��R��+��Km�ܽa<����B��6lC2t��a��8�w�o���9Q�84ꛣ����A5��I͖Q�y���&;��4ƑA�b���3�j��d��3K�uG�a_i����3��Z�b:�AM�mE�%�q���̌3��@C+&X����ɛ�9�>�>|� gyh��d�@tZW�e�F7�vg
�X��#%���6�er�d����I�$9(�+P��߳9�Jp�)������)C#�6'%������ZIv[B /Z6����:<���*�'CZѓ��o_Y���_��]���M̂�u�m�;�#�w�B�RA87���Ze���3ّZ�q�p,tQ�_䩮�-�]k�l��U�3o��sa�qq�U��Ӫ=��槥bf���*_��sb�+���ytt�V� ¨���uw7	�m"H� d�o"�JPX>R�L���i�'�_��v3��Z+-;�J���33H`��d�G��BYV�{���(T2�7DiK�+�ਤ�1|5r	�ĴUAK����O��"q������&)���@Cլi�,��-Ɇ�v�̊�6���VgKCz�Ɵ�1��7W/m4�\C�
�_�ݳ�<J�]�2恲�.��F#A5&e�B"@��\P&�0�5{��Ϡ�]<�jo��3��!N��*UR h�0��l��}P������g�.
�����)^�+�a?�ĩ���x/�k��-PA��1qӥ!~�)+�s�� !X�İp#S�<��=
�!'��&�l���n6z䪾1�,��G��]��A�Ҭ#��'�% G|��=���'��5b���5`t �ؒ�<p�bL Og.rL\��я�b��?l��o�zz��$�-zݿ&`F��r���AC7����z�<����#12��H����|�D��c1��K��q%WiH:}��gyD���w�B0J<�n����	y�}��w��{;	��CcA�k�z�����ƞtl��#hCg��檠"��&U�2z�.�Z�>�T
�S>��熛��C��+�������蘜�Cz�\�B�?#�E�#|)BLNF�,ꊤ�)Ҕs�g�A'�il*z��5r#��*�w�J"�2<�������	�A$�s�/!��L5�������G\���L]���|x�!C5W$����I�<%!�{t"��j	t�[g���V}��*,q
1g�H"���"�Ω��S%R�C۞�:b�n�L|Vc`q��&�>���(�M��r5~��"A~�ց�,�"�6�Z�E� x?Դ4}��1�x�$B]�|�zۊa�7M�q�Y�����o��J�r�%�☙l�f��7��`̨��C����~6�B���Y�"iX1���ԥDo�yJO�H�����^;��.i����ZܞJ����1�o�����@On��y�W�.lFL�r���%�R��u�@L:<���и���K䮺���lC�L���w� �7bc�l��T�ab�ÿy�\l��ſ�c\�1���,v[��,YWݼ4�_X�g��Z�L&w)���ߍ״n|3��KZ|�e;��J�(�\G�Sc߿"�U�/�6��x�}��̘�y�h���3K����?T���Æ��w��L� Rh�'H�Ͳ[|NSI����t1��H�3�r+V��4���"�A�=ʆ�b����7�LA����U? �պ��f�>O'e ��B�������aT���OS�6?�A�m����gZ��lAb����ݨ�},R��� ��^��R����������R�^f��.0�z�3�]q�O��L�*�]���.���u�E$��z�2���ݼ ��Q����܊��*�EF{)��V�M"
-���>�h��Wm�s=��,F�G��x�����7o�-mK��._�� �NNq+2Qih��������h�,�5�\\�ߞ�(Ú�,��f\����o�is5��0�L���g^\�O7����P�5��JǤ���q�>���;�C~Ijf�G�? ��/�Ny��_� MW�4���cmD�uMR�jFb)�Jn۪���p��٭H��dX���@�l�@��$�ECۜ)g��ڈ��z-��U�/w��5�P;��t���祺��Ga%$3pl��[���%�<�Si����6r�O�1�8Gpz<?d�a���E��	I���ۋ�=͟�5k��vOo�URP���UykׇBe��Z������f	��%�O�K�H�=��Z}�q��!���������~��
$���t��o����"��x����tE���ǥ�ELI1�?��T�l28�?�8@Ƈ��~`��ﾅ[ߙ0�M��	0��<��al�(�&��M��k��d4�A�K:Ms�%,��iQ\����z��&n]C����#]_�J⬾G���4�D��z=���d&#�F�Ђ���>uA� �����{�Y�~�?d�,m	cC|ҧI�14R����f��K���T]��� 6��
*� s���z����8�S�pQq���L����K�DP\-%V"�T��tJ��_`�Ä�)�-L�*��d%���CٖC��ձv]��4=�Pl�a�N�W~��(�'��)�-zsI��hKZS_iz��7�>b��E����H�=�0U����MY ���/'�:r�{�^jb��Րj����,����Fӑ�s?��h�� Vy?U��K�8��Im ��U~t �[�\<.JPVOn�8oZ��~�i^oB�j�
�ϕ�VB���DX��촕���5PcsJ�5; GS�g����0/X)pl�9m�F��*���f����e�S��}�Q�A��3�V���%��Q��S{b�멂�+\r�=��v[A�`3pէSn`u*��UVʸ���ӑ������V��X0��" ���z&Ьuq'D�?hC̵�S��X��(�@�Z~;�6����$Ɇ
@"IΝ� ��	P�Ѷ2��fy�!/
�����6	�����X�(����)D����V �LO(��fe:Fh&o��z���n�ͨ��Hc��g�����"S���ʟ�Z<Vv�~��-��f��0hI��t���ԯZ��z?�8*��[e?ҡWNacy���Q�f>Cs�ӕ����̣��B~a����~�n�I�O���\�a�F�Z�X�%��P��7�WʰxX�F���-P.)S��>m`\��4�f��kE|�q|�+��U�Q�ϹM%��D:憚�y��N�##��%8�;)���4�=p�^�(?g�5$�x�[�r��	��"V�}��gRs���W	�󎊷�hT�aPX���vv��umd�G9���}�de�T}����{�*
�VۢmV�x
���fM�ױ@�H���e��0ƛ�mJ���d����0�	mT�th5Z-P��@w�I�=(k�Ҁ���@�v�x76�*�v�'�X�G���A�dI����xx��M��W����ք;������\���[(J0QI=�knFL��X��p��c���S|��A�l�~���|O��d����A���:v&z�^�﵃Qn�f�ߨ��5�J/m�rt(��*�Bؿ�x� ҥ��4I�߈�@|^x����vS��	�bT�hѮ˂���n��=ֱ��\�3s���$��j� [�z��V<�*��.�����pT�2�yB̂l�����\ؙ[8��ld�n�c���U��gē�,�9�����d��XĩZȞ(ӕs�H\�_KS�U�d 2m�@�+�}혷�L%���]S%4ʥ���Z#��䳑t�\����"�}��&�a�e�hIy�D_P��E��&զ����r3O��tB��!�M��+r��T�é��������4<uЏeB��k[�2�Tx�T�<�"��Q�}�b0C�$�6���rM���}��e2i���6pǛ��$�}¼��
��<��Q�0��5��a [���N��a�"@?�wr�ڏ9L|��e%��}n�����u#�Blc��+�����)�w�²�-�R��k��V�����t�� ��Y�°n��̰"�v�`��4�[-r?"��ԣj�����S&�w>P�)wͤ�,_�G5�*�t��E�n�C�b�;)O����WC�u%A�8�*�y��ߝ��zv;�4nf�A2J��61
�؜�/��a^�.�G�3���&D��=���@�D�X���4�q윭ٍ�MW2O�7 ��*^���4�Y��Ù�y2�88�X�T�K�a�YB�������<tw�p�|!N+O����Լ�����|��[n����Z�c�;�+p��� �1@��{��t&�����YHᕜ1���q�Xx�/Ӫ��E	���[ri�]�s���W̦w�:Lym���~:�)��#`�aa}��<�1���+���$�8c7���u���N��ߤW����T�;�A����:�w壡��]��D�1�+&)�}\xzpQK�z�$����Z#�Ғ��S��[��"�E1 _̸�� %R� ���Y�I$��h��[���"����:�=����;���Fcy(쒂�tw����ɮ�_���w���o�s25�'��(Crxǻ�9@(k�x��hyr�K��kV���akMՂ���.�df6V�z0{;;fY����-;���xmہ@���J1�ǡ��������-в�J��M9u)���'ּQ	j�`��)����_S��Aܛ�?��܆� �wh=�����ДYH*������o��a"��!����VPS�j`��YE=E�N��kZ��D��aCH듖6n�:Ls4��cm�8q5���f
�ӏ�u�O8S?E����2>��b��:�YT�)���{	fKn��J��HD�0j2"q��F��k"xL��8�g���)�_��Q����}��|odD	Xx�*�lGuqt�(�znrz#� *��rؾ��V�h㪥���Q+��^�mp�ٱ��f���2�]D�oj��(bL�8*��l�BZ�KȖ���^Zx5D��K���� A��+K���(���=z�U1/���
}m|L����13�Ҏ<���Y*��ԨXI�/����F>^��[�K�!��h��n�۵�|��w����V�E��3�&s���KZ<Q���OǷ����I.�nI�͋��Z�%w�!�S�:��j7z�Lj(�݀a D6�B�Z���=��%Q
i���f�$8�ȃa�`�ul*��-0�WX�i�~�!Q7t����J�7��cWs:�����5wj�5�(�;���3�\xE�����ӎ�J�4����̒������c�O7N��C�QM��T.�T���~[�H�K$?u���H��ܚڦ>�۬e�Ңxq�:#nz��k�/��Z�K�S����� �@��&Oh$uCjN󳞖���8��
 Qk/��LAx3�ڽ�*g�ϥ�&�!�b��!6��#Lw��l.�r9�����h#�eOŻ)��N�ڈ~��|����kl�����Q�)OP�{����{e��DH���"��Z��;��z`����[������jlB�B=B-���:E��D+��o��:�c� �;l.����o�w��q����ƏX%*O����4�P���d.J��j����}�0� ����JUD�f�\D�
��= �7�dԆY�����:���ԆD�.54<�� �E��3_��9�^aF"�ž���av�&#n�+ ���	>QoN���0������,S�#����u����_V��V(R�rN���!���Q�9R��Y������������c��� �S	��G��%�1��m^����	ڼ�0��m�JN�)��-`Ţ�H�s��6ڦ�+�#�JO�i�� !h�߹�sT�����Pb~��?�\�Fm�y>w�6�h����Me�6���m��⠡�P�@"���{�M�~��*,W�ƨ���ʑ�4��Pc�#�'5���+?O����P�J����Z��Q/�T��e��`�9�O�f�IKn���9M����;%ק"��K ���Po��-t�_p
���Mx�{R��D�n0�^�!���I	���/�ނnu��0�|},�^�٪_X���C!4���ũ�Lwci�Q��Õ�<�l�l����&L�QdbQ��`�w�q*�UZHV��:��Y����i�jn̋*|U�gI�PmPoD��l[��q�8/��B�%龤K�,�|�������^��}�GUӸA��c�h�	+���I[]!�O���*��К�}�Å`��+��_A�D���T9D�2t���G����0��*e3��Pq8���KB��{� o��3�謠��Y}KD	զ���)\��tƶв@PyOc�x��:��Uk)�#PnG���R��v���6AiP�kQTZ��K�U��1d��,픤\<T��t��v. �A�@��+�:��W<�T�y/��U6H�| ���}Jݼ���7�X@��H���$�}s[#��f��jyoSѽy${B2V��튐���hqS=��NyN	[�G*���lܩ�	�-AM��ږ��U̢n��D�|e�l�cߴ�A���I��R��ʬ�"{�џx��?��Y��dyi����2� �^���Lz��2�g�O"OKj��Y�1��;�P�3a�Tn��Ft�}�M�f�vK�_�u�$:T2���s���\���bC��慒��jrh���:���~�M+ BtC[���--q�j��Z�Ch��;��b0��w����ܡغ|�	v�u�mb�i��.������Ň�	?+ۯ+2�H��%Z��N�Ѩ�ћ �p��"$➚����<�FO��e����Y*�A�r�f�"�Ⱦ4��r�!�KM�������?"�% m�r�����hQ1�ط�/�n��� �6+��:�q#R�HTgD��'����AV�ؙR�������X�u�^��$���?V�H��6A�Q�Jw���#�����XQ���%PS��᱂yAT�Qzա�O[&��#�`�y�X;��&����W/?��Ƿ_�%by�4ƕZ�������#{�je��J#���"���s({z���Ej;v��M��&�Y6�'oW)�M��l�G}���B?���_WI�<ѐ�� ��!w�1��E!�\4���l�� ��������3y�x붘*ӫ)�ȫ ��7��n�:�2��UE�A�݂�SZ`i��8	h]����7�~t?@a�MB��g �N��Sf���*��t�y o?Ĩ�(ℵk��Kt�Mfm�.�A�]M��kp5u�%�UN[�g��x4A�l���Ux��<�G��ꎱs0��+NP�u^v)1Ј�e��<*Ȝ��8:ą����H46�T7�x�Ҋ�M@:b�m�>�����qK��xύ_Q2��lE*�^��T����Qzqa�����Z�5����<�N�ߏ*Ʉ�[M���S�L=fZb�g��gx�� yȃ>'��m(Շ�j=��	᚞����y��O���7$
��.��f2��]7�|@�&�Eqq�d���k�v���y|BRM��:���t��?�úP�{���^�Z�^QU�n��uo���]c�K�r2���W
ʅ^]��̔�,�F0���6I���zM����Pg1�S��p��sC3��jZ�3?*H�lc�*�_�=�t���e��;o&�Q0_���@CY������KY�ח<��#�}���k��+޴��������i$I\!���,��%mi���Q�jsg+�YeіM(�ى��2o�|E�U�4��|���눽�|*�P<�uDW�ۃ�H�a�iqH� cõ���-�Nz�Pd�1w/����NBm6)�MBN��~���$�g�.,#�M��r�b��)��kɚ�N�bzD
=|��WâR~�bh��S�{��w!�e#n�B� m�����k��n���`@[ 3��i�!��J��������������yMwug�X�W�-�A��y���u;7A(8�[_ �T_˓A��I/��zZ�q�M	M��n T����(�W0BH)0�����xrW���W;?'X�9A�����_d2�N��/��sҭY�5m��� �J�ռ��I(�m��x��|��lէ�Up�)?�	�f�PW�����EP�nz�w���	 �
�&w�f�)��F�佹�d�O�A��i�/?2�4��$�l�y�����PC ��=1���ze���-�����NۡhW^��|��!�Aj:�G$��ӵA�H%�8 �Knb�������H�s6�/:@�9���`x����.p�%^��2��k~Y��zOdgɈ�_ Ii>hH-p̬`�^�=g-�k��� ���!�n��/���ϷY��Qё�0�WK)��1�q4q:#H���Q\#x���kf�|���{G�j�L�>����tլ
G���ك�x��F$|]&m7b������0��V��
m����c�����5���XI�2���ʵ��gƼ�s�}q�i�r���4�8�i�:>���G���\|lOຳ�� �q����ie�=�ݻ��vm��oDcM{�_-H��|&�wg���8�;��5Ԏ���P�D ����*����lL򓲩���#i���1Ҹ�G�;���D+�.��`����NH�:��Jܽ��_��hs[cc9|���	�VW\�~^̱� ��7��i�=?r�t�q�l��zF�3�v��1��p�<���ԉ�<����s�125�25ѹ&�|�|Y�)yaOmZ4���P���"1@��N�N)��J���]:������ch��� Ȗ�-&V�i�M���mܒ���Ƿ���*��M��T���B�{R}X'I�H���y �G�r�O�S2�
��=��ԫS;�No��.���	��꧆(y�:~ɶb;kr�eޮ�-����wy��~�H�z��0�ވtK0�-<م���z�����{ϑ�e��@�R�y�2Iz��؋~��E���1��}��wb��q�p����t���1��&2�֧4F'�W���ܘ�l��=�L��,K�BX�-���|Ĭ*�"�&z����g�|D���X߄P@2�����JqG��`�T�������M��jZ}z��Z�sӋ��	��-F�R�4�?lw;�$<*����Z�;�/.��9.P���x�%ݵ��`�ɝ֑dv����$��F��.���4���4:-�5YŔ$E�|9��|�N ��8���H��%<���|��q3#殻e��qc�<��Ll�K@�<�c�zzO�:B�g��H7�g�c��$F�ZE>F	�a�1�Qm�ޱ�ذ�V�����)���R�<?�ˑ�������( �_ ���.�b�o7, }D��4[U4�˹������(a�
2:�5xk*�R<<XUP&��!����q�6kdP|��U��=�zZL�[�OE
����x�V�I��n�)Ҝ���M�SJ�#靺����.q�eYo��ck&t�!��e.�ɰͅ���9/���$��n�d�B������թy��T~��G�-�忱b� �A������_��jO`6�PUu	�"I�T1�!%Ճ�>����Ko��8��Om��)1�L���8[G�� a�9g���?)��=}`��X-�*�Ϩ�u���Bd ��`c��]f���@^b�Ȅɿ����go���-�9䉥�<!���mp�W��<8�b�=q$������� ^���@�:�6e�:�b���+,��h�z��,�j�z�"����Q��x��l���Y��
�R�.����	,����>�1��������O��P�j>��J�p!��h�����/cx�iy�&С(�8�l∊o�=�����g�T&Q�C^{ֶ.�}���.G��-���!`AS��(b?������ƹ��J��T���e��uP�#��jA����/D1T=�;�\�� ��3o`G}� *g�ص�{�s�jT�T�j�rJ�x�����C�S銛�	�Ԝ��s�*fġa��`���5������ǘ�VRp��]�C$�u�,H��6��΢���Ied^���9b�pu��p�B��ر���.c�%9�0�xے }Փ�I�i��|���ܴ�ݦ�Xm3k���Bvz�[�Z�3�ޚ2�Wo���X�ݑ��y�9����������'���u^�g�-j2�ԕfν�m�Z����Ef�@W�t9��N-2g�{@�l5,$��Μq)�-9<����v"�II.�|׼��`SZ�<fPH����[fO�k�`)Uz����&jW7~�B�qB��m1��a��6��3ɣ��NB"�D.�=�|#K.H&��F���i�YK(I*$$3'�1���,Ѣ���H��wUЌ���Ҵ���( �e/�@���E���|��
��F��8ٶ1��������Πz�31�`�[XL���&�F��'#�l���HJ��u�{w��������������J�*[�c�Q����зU���#L�{FSڦ��[�k�3��Ra��d�^�^7���{��
V��6u�6U��Nde��H:;
e���ȭ�����N�c<!<�뭶��R���A/p��l�yz�/����8�F-de��Y�3���%ԣ�HOd-D �Q-ͼ�!�t��'�����ϯh�:�����p��4��7�e�W^���� �b���T'�j�m:HRK0Rrvf�EFK�n*��f��R��'@�asے�،�(^W�Ŗ �3%�@��/!�?�����A�ΐi=;P������&���Qš�r����ȌH�׌S9i��yW��7�^-��R��1omv쥒�i����a�P����J�h�ug�tH�6�=�EV5��EVu<X�π8O�e������n��B��p�Ψ�!�#&n����sSC��m @/΁���g@�h����1��N;��С79h:��0Z���|��m�i�I��P	$8�{�?���>�Ml�<G���_�M���Hj�?�|Ͽ��v��7��H4в�eX�_D�~��ǚQW"��!!� ��P��������΅��@ɭ?^����LC���=r���:���9����}����<�/�����H$�t��QTG܎hٚ4�L�2���!�Ej�9��b�dS��!�O��C��AU���8�����`~'1�A�<x܉1&W�Ӫ�/|uj5r����o[�Ċu��E���i j��^�2�q��7(��Y�����7���&����$Cw��7����N�U�ş򧮞�jUrX��>H���Y&J'��:\o���\�3��ɚ*�t��2�|,ƙ%��c��=�a�;�ס)�(�u�/x6�iQ���C0�`����lZ&����&W��7�C(k�����ېa�N��ܖ6c�V�
�<���)E��m��D��zr�մC�@F���4��w$ۻ�ʿ�ΓK"��������y�Z\�Y�딭j�F�,�h�ֽ==h#�2��U�Ʉ?(���>�Ä=�6�r*/d��
S�a��v�0�z�,!�P;���[�R�_�2�X�X;o<��0�4z�G6��������.�6\����.������G�4��s��xƏ��=񫡞����4ɄU�2�	9䈑�������in��2���WC�>v=1z��[�Z#�I���HP�b5ƨn�-���P��T�/Db�m�i-Ĵ����Uq�ky�L- ],c�9:�hx�DL���]T��y���DRUo���K@�W����l�"�sx��G�8�l�9��CW������oʟ�e9g�p��Ҝ˸b,f� *��F�3���Ee����H��0�� I��+�On�ܾ��_��6e��,�|���&T���J�934�~�U}.��1���h��mӇ��㬔{��BAW�*�����V�鸜�%����X��A*�>�m���-�U7�ѡ�t�k�tԑ�U�Jc���9͉)�e�$O�C6I_�6kԌ�Dv=A5�.�L��ݓF��v}������^{���I�]�z\�?�A��^EU�H�4��l�ض:~��_�7G>��2DL�3 $��ϯQ�����]H�(�d��/�g#��]��}h���}a!۵ۙMKr�:X:�l(d`��Z�a��W�V ��@};��
���Л �PwH�±<0d�����\s'�7��V O��aZ�������9����q�0DR�%QM�,���1��؆��m:��P�q���;}O�#��~��@���;�vx�	�l�j�~��.�ޠ��}�X�@ �eP���N)�o�N8�eDdj�R�zG�:��Mɰ���j��;*\�o�1�hS��d��o3�O/a�KxDZ�-�$p�1/��8y^�!&��Ztr�z£��e�}�"����.O٠���)ښq���.n��T���\:>㥵���\�cBѩf�����p}�����D#��%�"ѣ��5��S[����/r��� ��s���fo�U{=>�
�͹<cYV27�w���MY�c��w<�'�u�㡼Q���-D�u|Ɵ̋�?�A�a앰�p?���L?��V
h�yc\dn�k��%��R:��=�!���wf�RP���V	��.�7?�� ���������8M��Wދؘ�@���pb�\�a���@ݟ8ܤ�e�o8���	%6��L#[�uG&��:���Q�mP%���h�EJ��V�>nQq�ۊ�||�X�ޞ��'c��ov�( _^-�ë �l^�9���HyQN/6�C��W��n��?�"���k�N��YH
y��V��k��RՋ_���F�!�
3�9�y�bJb�ÿm#~�ڽh����>�*�1�.j^��cw�c�r�G�iV������#�]�'�K��8�;�{���W1�Oj��xq2ol2.5��n�u�}��3�5������O�Z0�4�z�a�b��ӡ㿃�� �]?��9���D�rb[FO�6la^f�����=�и��_��H�a�`K��8D
��@��幅�]R�`9��o����Ϡ����}���Ǚ�%�!d�o9	�,AX���U5�i��|Jx�\�9D�l.埯�%(=<��q���h�~0���6^�⭌��^�EIi煕-�����$� S�2�/����
�iq�Y�I��	�����6�_S�V���ꋺl-ݫ�����`F��T�LE�'Qs6:H06�GP�4��K�O��!4�B���v�Pϡ��#���ۀ� j�h���*4�*�γ����x�<�����9E>����y�{
@�x�2wij��o��q��~���2������,gl(ڻ$�hk����j��unm(Xs�)�8�>>Dy��~� w�>�)�&�T��:
5l�+/���k	� ` �`!�<Ͻ���^Ju��28��^�$ML�񅾻��'F���t����!���W�'</��|RƋ�J�,6�\J���`�,B��D��j��&���A��zк�]y�,����A�u0)<Dt�u�]��n�����%�{����,m�A����IQ�6~�g���5��Y/Q�r-�6��p��E!�$(�׉�q4c$*��*�Ir�î��)y����-~����Xf8Xa���@ �̔K	@���i����Dr���~�8��� }�� eɩ��-^� �{��S��� |�<W#��Hi�Ϝ�<�d>�O$?�͏^t�fg��0&ß52;x�贝�w��~c�㬫okw�-c$�.��P�b�JDd�q�/��qKW�22��./�1�j@>1���]Î�X'!j�N�u��- �?#9��8��io0�\�3���ul�,�\^�\��Y�&Ct� �,����(D]+��&#% 2�(���u�V��;V��B4h�W���2?{��L�`9U=O���sB?����6�_nf@��`햐8����0�����Zvf�(6�#p�E�Fpgǌ=��*�zjU�G��=�==�����o	]i��Iq��|�R"��D���l0B5>a��S�^��&Qc*��Y��+��|lMe~�^��V�lK��l��m*��}��I��;Z�	�؀<��P�K	(��m
��B��%|7O@��M���������G���(��(%4��A�'�e�#�8)��_O�����>���`?��k���e����M�*��.A]O?:�)�YI�,�qm��ӾH�C	ubǖ�J=���J�<&�/� n�}y�Z�l�����A�cKbc��\������䇙�<M�HxYޱ�,��E��DsR�z��C5�>=폙��5�Ga������Q�9/�]n6ŀL�)g˴AB���5:h�6
�N�2{�eA�1�~.�k<�r�%s˂5���5�#K�e��nwu�)�	}ޢ3Xz�G��3�S)�]�;�p���96�ct��d_�/;2�Tʵ	���z6�:'��;B3P Ĉ����v{OLm�����d-���	)
U�̃tmᜨiB�z����c��T�6DH	�;#ƸXL"9D�/L�J�	�J�<���'�'���í��ʿ+�[V��w?�@,��c��t�dK7�eX@7в�r^�#�8m��-È���ѿ�A�"yp�T�C��GJ�T�gY�4�s��uV���9�,fTz#�}|��	�ڪ���	����&d4j�&���; &�)��򟖠D#��ϸ������'E��B��>G��%u���L��zJ��_���Z��5�r%����p�ne���������<u�Y�?����%���6FS���|<w<B��o�O��]�afǤ���=9�\��1KʷFQ 2����ɶw��l��P6:�"���"�I��mp��0�W!�ι�k���6W�.ˮ-��*�/HE�
 �_0����8���rT �&�@�j�*q��+ܕ��2��!%%�Ԙ{#v�0��A�P���dA�e���0-�b}"��R���(���;�X�����4�Z�уy
1��-���p��+�6����k��O����Aq2v5�7`��dI������j��g��/���JiV/sC�����>9w��6��*=QG����,א��.�5�'ܩ��'��7a�c~�oIs�8kc���\3��`{ ������=Z)����`�a0��Y�3�S[����,�5� �]O�rl-c�õmE��<��;c_�����CPAct��"Q5MEڷ���_4ITw�D��=�va�2�׬���y�l���<�p�HV��fkd�5�d$��w^�Rl"R�ґڑ������	À�_���=�Ɩjd������
'D"���^^X�����u�r��Me��E���6�0wH�'\{g؃�V�`	F�6�g��|�'�#f�\| yur�"�X7ݙ�wJK��Χ9w�_2���.����l��X'����ȫ��,bL�����.��پ�'6��h��� ��p���3f��W����'�IL�9���ĺ��KU����N_ �D���1��mþ�}�Z߈G5)B��4B�6����Z	"w��ϯ�%��5���s�+8�NU�����z�2A�]�P�0��p�������=�k�^:��,��\a�ś�gs��mw��V+Sl-�y��g�*m��ű��l�Jq3y!;=�`�c��梨�&���������S����w�m�-�0]�N,D��%L���oy �=5��G܎~Yk(w�n�C&oO�V��ͽp{t]��|����d5�0�6�� �<������Z�AxuX� Z+�W�2������SrU�$�q��������ܼs�U��k��Oď���m%
��S/�A���/�wk�F���7�`蠕~���E/�_ �e��F��ڏoy��e��x���P�NE��]���=6�͗nf;�9�y�>�g��^�@���N�������-�>:T�@�ɲ��C8�'Jδ��Ý�^QՉ�l��e��z���>��}�UX�k=�8ƫP/Z���!�O�2��o��U)��Fz������O��8V�XM�$�6e�ƴ�jc��V��R��m1��E;3�c��R�q�趚���85�6I�f|���������KW������^���^:�?�n_a0��ۘ��q�$-Y�%�� ��x������h�M���"'~�����MQ��i�vO|X�й(�ermd�����#U,%�H�ݘaFn�Oc��ˈ�vu�d�����r$�zsq��ǋ�_��˓�ɀW�bg1A�¡�V�.D|�56���K�Pd�YW͌��#�1q��?�9e&P�.
�zY"�������%eY �		|a�m2�Ch˒��E5sy�9�*��Cy���E���-�����s��vBY�?�9����ay�U}Ñ� �l�ϗ�.�cYac�N ��p q��f�㹁�Z���������Q��)�)A��S�W;K(�#<[���]R��%�?�%>hP�F��^�H�413 ��WX[RkK�վx)��� O�y�ö�r�ͻ�hX��yL�i����3�ހs�?r��l���3��뻺Ggp��`I�l��[?�n�G��&�<�fP��ۥ)�&{;R8H�E����V}�ٔAi�����U؞.�l�@��������k��RM� A�wg�V�Tv#ԫS��Jf}Yt)΁�A�"8X�J�`�&yJCf�����wN����G�i�R�fy����Z`�������<�C�}���3 X �e9I�P�W�!���N�l�&z�W���-:�4
c�h`�h�R����G��T�C��3��ɠbd�| �iG_�P�:	�Y�^[��s�5Ԟel��wV�W�f�2g��Rr'v��G�6���q�r�jk�u1�Wܵ���(>�i|��������"��ʙ���|đ�K�d_ց�م��qsL��q�*ղ�H&�!]%H�N�c#���i.��dZ�Ğ�L��$ngY?����V��� >k�@�|T���a(�&$��j��f[�@LH��x2$[��D��A�Ȼw.�"�u�X�.o%���.��-�XPv�O(ϙ{�I<��4������px�r�;�e�ǡ(��Q'_���7<ㄪ1�6�wFh�_��Շ��)0��:l�B�����,珳�#V��f �It�d�Q��W<L�Z�EA��w�Y4��`�F�!�����]��c&+z�ݑ����
�&�Q\��fe\Uʅ�0dǼ��Z�7�7O9�-� ��R�V���Q�m�7t���hM_��hm'��ʁ��}�4�L�A���l3bJs�G�kղ�%�4'Dܷ�BWi�}v��yV��]�=xq�4B����۠�YW�b�%,�f�s+K���E(5+%��UP�.KU����Ch�f�!���&R����7\.�Q��V����@��Xvv���������%�|�m�]�O���,:.w�aĵ��Nz�}�	�.Ԙد\uӽ[�b
F!� �!kl�<gE_��/�ԛEo�����)�ɝ!���0�����>��V�ͤ�������rۢ�2l�4a���x+���)c?}N���G�p�z��(v��e��ʷ�73���s�y��>I6	�+�/ �����o�P
�iG�eh��B�ID}"<=H^���c�8�������n��
��)�ގ;45��C:,��ns�Q'�B�S�:�7����:{M��	)�+������w�=����88�ގ����Ԟ�+�1	��a�����Q�Ɋ�r����a�1P��U����p��Ը�$s�VԲ��]�p�>g��z�]@˖6i��'kM;�24g�=b���N��,p��7�U@��	+a�>qN��=ap��)v������ժI�r��c�P��,/Ki���"!ei��-hZ�Û�x!�?�OH9$�/������ԍD��3CA�g��t�\���CiÌ���]<�ek�MCV�-SĴ�h�f���eى����ߕ#4���0����ָg2��.BW~�&1a,봈I�x����*:���C�V�"�r����d�~x�-#����)����K��
B�ЅUZm��>���e�z��Cn�,,1�
�)�L)&�� �O-Ժ�/��L��u9���U*?%�Y/BN��ʰ=nn�i��B�`�T|Zn(*{|b�nwJa�ߊ��*���	26"��I����{B{�E�
��~��v�(!�V�X��w����Y��������
	�|Й�]�M�h4����&�����^��hR����;p���^Q_���lE�D[:6���}e��Itmc�}KzB"B<!���Z�̐��4EN���-��x�f�Xn?�6'X	��'ح%�C���K�5g�S��zcg�pS�0�P�X��Ie����0
d�u~����o�������>>͉�����	Y~�u���]�9I��p���2F�VM~Ab�0n�C=�J ����cW�
��Lf��ʥ(\h����S�Cb�x�kleO� ���W҄_?����?��PG�2Гݵf�ഋL���Vx�P���s�JѦ	#�v/�O�e�$��L�԰pn�!��h@�u�1+5n�Ad�єkS!�	M�0;#i�k�W����7���J:�iLT�
Tr����8̈��ձ+�'�l�Y�6W�H`5�V_-� ��ef?-(�yȯ�w_s�_:g N��n�TXƴ�9�j����LWpꅆy�/r�����0���T�)Us�(��à�ۑ�HxWt @�֜Y=���hd���b�`~[�M.���J�EE_�,ɠ�C���"*�9?�H�p4v�QF����R��כt�;32Ҹ#:/n+bNM\F��o�#k��F�r�Er8b<jv׊�i-��Mnco�Q��������:�LВ�w�H''�����c���RË_NZe�������Ƒ�E�jB@�ƉgB�6)�,/;!
�c.�j�B�%���s��;��mj(g�:(eP��͕�ێ��o�}��oR�-�$���Do�{��1j�j�C�:;���Q��%��"�g�I��l��U�7��nZ^�ß{��_ۖ|ݢm<p������7��F��O7H���YТN��jaa�U��Zӯ!4�Z1��)	��?ي��|��J�x���KS"���/F�mm���4T)aZ��So����\������1ʦ]�n1�z%�wb��!y�n�����0ZO��<v{|`W�{��`��[G���6����W����1(�S������f��k�e;Aɲ~�c&MǭJA��\{oG�K�ߕ�&5eYq�$�;9��LL��YMՈ�Ix
{ |��� ޼�r'��:���NZ)���ʢý������[���?��nڴ�eV��Y�	ՈuWN%NIG�^:&|����@i��\4�u�*�%k=F��]>Y�-~��',[�^����T�+k�m���EU����)w��NBpŮ��M�{Ȅ¦�(�e�C��b�wuF'����90Q���1��P�t��Lkݴ�["Ss���1�D����~��~��j$H ��'�Bf���L&㑾��~�*�h.�u��"3@��g �d��diHu�u�R=���0��V�W፹�?k=�sԋz��]����΁��0nl`�?T���D2������^4�^��T��Pf��E_
�F/�̱�����zZ��4�4��4,R][��iGM��?c�%b�;�p� �0�fپ����fo<��S8��'Ḟ'��p�t�!*�֊���A,����2@Yt��9�Qeݥ�+h�@\��t�m�鼋:'�rn��ӯ�<���veI'�2@�#���6�
n7�rƾ!�
��~�l1>It�/lU�x�����T��}��Q�lτdb��*�Y�|���.=�c��U�?��_-�!�k��h���۾��:T��]�Q;A
x��ϖIb���f��V27���'`�����t�A���-p:3Xfi�+����}����2%-�L�U���˱���oG	Z�����O�o
���=c��������F�� �,��t%@G�Mݯ�˳Z樜0$�Vg�us�{E�¹�%��:oZ��'�C\E�ce�H7������S�}�����_ì� ��S|l��8"\2��ꒈLa�6\�[��� �)y5���>E�m��+d����}[��p��Q}i}@Gg�4rz��FCe�r᫓w�Y����\����WG��:�������Q��|t�΂"�dg��Sˠ�O��ނ}�-L�GB;(� �b���@<Y�HSA�:�rr%��q�	#��Az�?���_�����8~�}?�[麨�OG���݁���P0��A�1����z/�p�HlKVkS\��F�n�5�N�����.�P��ۨ��#��v�j���v5�"����oĴ'L�E�5^�{m�*�٣v�pn����t����>�֕B��(8Q��?���r��!R�:�c����~����~N�qW�d���ɅD���L��a�������s~��J�����@�0�,�i�T�aW�Vr����kO�,z���"y�Q�x�H�,�P�(�t$�ֹ#8�&ҾB��2���`�7s��}(Ӱ>m�T� SU�`/�h.5LS�2:�������P�~&2Zy�@f37A�XjI�[��|�9h/���a���W���rT74(#���$Ag���a�2A�R�ox�[uF�7a�.������2�4?�t�z�ۣ�#����WT�+w�o�Du��\*̦���m\��]ޒ'��b�#�X9�Y��Sm���sPK���+�(��L5P���.6S���񩉦M�P���eN�V�o�+���O���mvP�f��%FL�T~�߀/�v�xJ��,���Z�{�)��K=��Y�-[�È���^��/�f����x��P'1���(�x�ӪS]���G'�d"m�ɲ%���� �/0��\Rlp#�"P8�B��'@�
?�jo�w�l�s��]���ss�����cr�b���������2��0���F�&�1�T߀*%�ë���$Sƪ4���W���K�V�V��$���L�k��_")����GM�=���S��2Y�w�u
�:�g�IN��~���g��s��Y-�-�ԾZu����#*�W
�:;�O�����H�rSG5���Ĳ�8�y_Y��ݮ�������V;|:g,��^�Q�fϥlϯ�Sg��"���C���}�\�\9��=�f�ç߱YK>g?���f����!B��[�hŴ�l�� �,_Y�Ӂ*�DA��9�:BRN��vi4~�$[\������u\�׃=C�%�ۻ�q�w�M�|o�O��3Q�1�dv�f�<Ŝ��<`J؜����j?�}WO�0ƒ �R@��������9Lף�Ht")zP�n�� i�)�nk�\|�����*�k����-!Q/��N� 1�&RN��{s��g�+VP%�~�ģ}��}�b6���xg��wP�J�.=bV�lĚm�شv��䇬h�
�������j%�����j�^�*��H�S7y��@����Z��)!=+�IP���2��[�c�'�� Ŏ��գkm����G���,V#9��{��q���L����! ա�i>R_'����;K/�7o��{ݴ��3(�P��c�Ak�J�)*��{�c�`���{8���g�y�9�$. \�L:;z��T��Z��r����3W����ȍ��I.�qL�5l$J�^ܚ���ݥ.k.O�:���4ڰ��2CLܴ#�"Z��j��6��=�蟯��"�Jّ��v��+��e���F�u$���������Bu��z�Vu��b�b��O3���=�E���Ʒl�t״X"ɪ��E�F�X��4ω�QC���5E�B3tWc�ݶP�4��k�(�M��B"�#>�+e���ʘ�u�xL��3$"�������f���+x���--���dx#���⧃���G�}M�A �['g=��
��%�����i��~q=2��lWrFT_)?N�w�,đ�݇�a JY�fi�͘+��5�-��>n�ZS8�²�V0�x?��x�e,�|ڮ�<�P�"t�ȡR"8t0�O�]��7�e���+��*��QV��5�R�d5�{�3����I�D��� �	/̭�JB)���Rx#��4dݝ/i��5�)�8�/ĳ���Y^b!�����k����8��� ��`(Xc���$���G3��Θ�R.;�y���t�Ӝ�Rt�T��vڹŠ;��+�Qӊ��M�!Y)i�Gs���x4��pV�f=�����٣A�v��tfH-��/�G���F����:tֲ�8�f{�پXV�+����[Cy[Ep*�$�����%��Sj)���cs-ٻQ('���f=9�8B�LtnWbk ��1�2��Y/Յ���q{��xh��""@� �OAw��ni� �|�~�΃��N�� F ��(���i� Tn|��sK�^�����"�̴����[��3i���5G��XӔ�6�l�%%��۟�r����h�tnP�����F���o)
y�ѿGOl����?8d�s��-��N2"��g'F;�^�`$���V�R�]:�ҥM��;CV��~çaQ�G	�`��C\㪓3�~�PҞ���煖mD���?R#�]�P�CgZ��~ʕ�[��]��è�J��kq����w��j���]{�l���\I�\L�"*��z�%q5Q��/�=�	դv\'<, �@����_%�ib�+wT_�V~X{=R�N�Q��p��L�߉��zL��M���@|�d���$qW!�C���6|�~�<��}���ӕ�2�-!;��t!����kgq�� c��X�4	�h2�mL3|d́D"�P�R�g�c��k��!}�V-�����c��j֘����);�~�"���L�P�	qQN����V%��c��*�xSh���w]�Ο}F�h#Ͻ���5�-Y��1vD����Fԯ$�?�m�l�[�bhx�@�#6(13$�du����:,$
i�6}˘�q�Ɠu���!�!�B
͊ ���^:L�Љ�y<V�����[��r����^�w�p.��o�c�o�?��8�O�m����(�Ѣ�x��Q�\�s�F�jv"�҉<^��?
�~Jצ]�4�~J%4�����Qԓ\�P�r|#h�5��!��t�<7���'��j뻆F��A�t�R��Dy�,�6�_�7I�$�(�y);�U���p����%������|����۰�Ŧ@����\%s�����r�6BN8�n�'�P�U��m�
%�+r�Pp���IS
���dT���l���i{���F4K%U˶��0��φD5�á���v�2q������8��~zz�Д�*�b�����pj�zKʅ�")0�lZ!h��][��KN�/6M������χmoI���i}��7NxNP{�@>-�R����h�O����>����n��D>)~��&��NW�:>�sl�I/�!�z�31�<,[{|+3`��<������Х�'����Z�1�}[m��U��nܐ��%
� ���F��n9ie�g`��um��췡�[a�W/}���o�KN�v�H�C��5EwөT�sЀ(�Y�I���ֺ����k�Dߐ�8�D�}ݠ5^
�Q�a�	�K@�d�����:C��Z��J��o��@-�!���aSgE� :���'�^�4�<���z�%@��(Q��I1�\�Ľ�������2�z|��f?�����pk�J[θmp;�cov�� �+���;�d�x7��j� ��`� ����c���:e����K�j]�x�>R����E}�thȟ�����twH=lAI�$�n`~/���'���C��v�c�d8��&����H쳐=��ڃxĘ=�x�آ�BY��y��o�2���>��� ���<��n�G�q�c�$��{$�3}X�!b�	,x���f���*��[i�=�o�[�9~�w���){X���>����s�IЇ�K^%$Z�j�L5�62����r�ε#����B�}-ܿ�x�m���
��yp�2�o�x�<�b����L_WK�Ӵ� ����E��lՓ��M5��^���ĕ%�`������H3�p��.6��Y��ȧ*�pi��@7$h��*��Kc}�TP<��-c�ᗫiI�92�kf�� 2���w����]~( ��u��;���yg�|�ZP���&��a$Ə&���ۡY�4��8�Z���y�c�~0�kח��؏f=�8�jq(�"�D��Ֆu�����̛��콪�XEm6�	D��n颟�;�2�T�1�/d!m�n�2S.��vf뾲�fײI��)1���V}��Z]�ζگH&bv�iq��U����l����giLQ�rǈ
h��Ρ M`�FJզdG 'a}1*�����24\�汷|���c<�	Ȕjf{H%�?Dx�1Q3C�=R��}X�V@� �ʂ1br�wK��w`�F+�����S��y���
�������D��uɤ�.��*6��3lYC�p�J��I3j_lu���F> ���i�]!��V]���%����O��1��K�O���W/s���-�`��U�K�A:�,�X���w݇� �����=׊Ta�Zm���_c��m���"�I(7-\=r䵛�!ثl��n���Ζp���H�X!��1����A۷ύ��7�~vЫ�um��=-C�U2��}K��%���B�	�L2�oQ���VE*-e����.����,�I+��m�6��17�y�G��� 	( ڧ������CB$x,�}ׂiNQ�	����V�?�Q����xQ:ج�E��)v�j��:���K��^���DNʏb���m���ul{�
�ͭ��pu��������[�~�Ql8�6�]݁h.f�H��(��j�ַvӄ�=#��cB��U�u��Ʀ��a�YH��	�6�m����v:B&y���i��j�I��`��~��wFֺ�%4��YD�7O�ν3Gm���� ��%�C�H�o�X�P� �s��tA��t�\{���=Ț�U=���Ϫ9�?���^ �T�����O���faڎFWP�\��Ͻ�b�"/�^�r�F�Ŏ��&9U3�31�2z�i���*��.ƾ���: ���Ao�S9�/��t��\_���4>֙-���f���ah�����R�.@�7Yj��TҖ��b9@\P<�?M�QO���kiY#�}=
�Mk5,0��~�yㅰ���]�Ek/1���hd. ۸�smZ����^ui��D��2��R�L���s6b����,�o�6�N\螓��1d��c�����h���h :ģ8PS;��v���b��f���|��\�c�h�]i>Mb���U���d�I��BN����M�}>��T�:uJ��� ʍ���MC�J��*��UW�f�[ �n!��h${9��GNVZA=9�4Q�-��)��U�+H-�;���P焾峘)@����\�_,^ü�U��1�,��e;�.�C�[U%��l!�Q�0�i0Hۨ�ҹFQ��?ʦ[��Q���>}�XH��wlG�ŷ��>^�p䙳r��	�")ؑ��������J��<w����9��rK��Voh��+�)�2=ݥ��Cm<�Vy$3D�A�9Ўt�i��W�Z�X�4������&G�OmUE�J)�G�R�'�� �Hqbm'�`NH�aڴ&�7Q����D�3��KF�^��p��� ��X��ThȄS�ĩ�����^G���O��5�X$���J���7�d7mQ�w:*YٽL����,�T���{��r�d5����R���\T��DQB��?��@��q<���?���gAQ��Oەję$o������\��HYj���ls�VF�'t�|Z���3Hhd|�F�@o8��ˡ�FH �x�Xb:��b��W�:�7��6�M���7�x�݊��T�ˉ����"i�6`X7C��QH�Q��e�y'u���P��w�1�zr�o�b�1!�,$Ø�-�fI��B�U_H�3�Zе�BǓu�2�q�q�qq�߲�%(�SW6;4x��Z�@� *�{I���qվ5W���A^F6>{��'.F�K�2��k����Q���p�^kx�KJ� ��p9#,�zKx���{�v�ymKI�<J4��	���m�� �2h�b�&�U�
?#�ݬ����Y�b��Y�p}��Z}���~����2	d�ZM�տ��$=x�`↚�:^_�	����e�+ �c��`���E���=P?�5�Aƣ�����6��Oy�].���ע�F<VM�˂/_���(���W�wM�^�]ǉ�`����3��[A��泷}4�`�z��w7F��E�F�zc��m�6���
�(W��QG�pF�?�T����j�L��T*�oc��LP��~����H�s'E�Yv���^����(;YqU�^i@�C�qkB�(�IZ,Uy0rE��}-�G��3b#�y��ܗ��x���KY0��S"��:T
k��Ncp��	��9 �䭏��hۂ���٦�;�e�1>~D�G��~GB���ZJձ��� D�l�.�0�_[�jJ8�!�kn�NdEe���N>�U����53Lz��2�ȹP�N�f-6b[�rONtؖ%��p������g�R�7Z*�б���^9��ȿ�
$N1"����%�Qo�˙� �vh���KH�ʃKȔ��xvK�)�����q���Ļ�o^�<� �f��x?�Wc�9}�y�a�t��;�0}���*�i��֛!��^���R=}/���zR�A��o���(x�˰�d0�R2�s�ݣ��'���sA�`�i��䚃�rm��a��D���N�w��A(ت�kH�PQ�՝��"S�"�M9{3aqI�k}9��>����=��Ks=������[�mk2so��[��x*
��R]��+U\P��0@��sY����fi��@H�����X����;p(��'�L6a_) ����G�T�0���P��/(���Np,2�&�~�QI[G
G��Q�T+�S���b���{�7I2��z�z��\FP���\i	����P�2����`�"R��Ȭ�xm�XHZ��ʒ_��wz����\�f7R�n��D�;��I9�C�aC{~zXE�
 nD��eN��)��H���9�&d��x�?k�Tm���Fr�QƫM�|� ��eOd�cFU�^��j�wf�@D��o��Rc6s�@�ju�e��6�xǸ��mVf�Fyo`	+�_}X���h�T�动�pA��J�׍+����QG�d���O�wMn<�\ϻ���\���%�R1��Ha�[m�F�D�ث����a�C��k�'�ml�N��:�u}��*�h��S���VP�aH�(*aݰlA"�ͩ���j��%��$oL}���LR��x5(puE��2��`��ܤ��7��-p�!���|1�C����zSoW���(:��ͦ�L��C�������=��}�`��_VGߕ�,��6�?5�ٳ,�^˺:4�HdΧ���V�/�R���D��=�Ȣt�������3���%�-#L��N��si%W��|�6�e��\'R����vX�V�VUlf���j��Ժ�[�����D���b!Tɱ�{��$����P�AkiaiG�״&\���Hp:ܮ�8ҵߵ�c\ԺF0{b[���l���7��aǫ^�z�v\�.���m�e�q3�:I�;m21wT5+���8�.d�e:�\_�u�[�P����+M���+\uh�C �t�5~��-W���i��6u�59�(6��d����{-.*�w%ࣇ�N�`H����kX�}�j��[��O_�=qa��P#	�
D�u�/�5&��hzF�.7���<ig��p?z�ΏӸT�>բ�;&rt�c6�I��v��æ=�I5@�_r��Xylw0���}���&|���\T�P�5�7���UA����H�&O�v��U�Ʊ�y���o�6�?G>L�3�d=���I�	]<�u��(����kzW�%.�̱��^����zX F(i��Q���7[�����!"�,�p5�e#m����\tN1���%�<�U;�[(M,)�VVgs ��n�lŮ�B*E�CU�I:Jr�N�׳A>Ս$ZT�h�w��o�� �!�$�������9٧۔|)��ѴtW
�e_���d:p�̛�� r���V��Oa�K]j��s�Xk�8<6�U/;�f8��^�n��Y��k�a����kOs�$Q#��%ӟ��<�S��$s�~���12�����	а써�{ns'W�Lɳ��S@
��H\1)m�c���$���/���bL��۬�a�x�eZ�C �tκ�JI'��=�W�X�9�-X��C:��o��\��[F'^��q�$��l(M>��mE�i�������k�F���q�ӺU�c�@���������z���3��^nHg�3{>���D�|t����UgO̵s��K���*��ՅO�n����5:��2������q��F���-q-��H�}�ő}��`cmseD^� \�p�W��p������+�B���������ݵj�6:�>GըŖ7c4��8��6�d1.]�yW�-�M[F$|ݦ��;�m�G�0�~rW��W�DE`VE�����,�R��1q�|<�U�%�ƫ Y�AX涌ɝ����/O��3i6�	]���h�{!���*J�"�ŉ9����J��?eA�}{Iv���{W�U�H��M4"���Dy���S �u�<Ӑ�� I��u0"�-���VZ����J���G�9�]�V�߾�<(����AwX�F��]��Z戭��//&7��!���>0B�,�ZC��X" �׹~�����o��3��>�Tk�L`�E��m��yk�ճ�U��Q��N���c��buV���&�������o����vn�����j�;����������n��{e���� ��Bi�����,��
v�DM�M��;�tF�O5�q�M ��t���u��^��ౠ�gw� ==�	�Eq�[�Wys��'=��#t+��c9�q;������պW�0��z��	R|����
-��`�����=5-�#� ׽"y}���^&K;�!�V�L�7�P`D�����B���%�9J��$`g��0s���	�K�����Ý@��7��*>s�
�2~�
i�o���UdUe!"�C�)	��`Ӑe��hn(>B�'�.�XL���+�K/���e�<,��IET�G�I�����<bF�
O#��%02F듇�<y�Ry#l�L��Lf�0�PJ���b!�����W���ϕ��>����� 붓�wH ��͇ۅ�m�bgwc�5n�V�9�k`��q=�Y�5+,u[H�vӜ�!kV�Fjs����I�����7j?(�ͣ�+�)�y�#��o'�붣r�lT�x�ߢ/�FL�h�zI�4n�_�6³��IF��:��)g��$��unE�l�Ƙ7;
��E�j&f��0�+�Ǻ�!ԁ}p�l*݌Z]4~���,8�D�A���a*����=�`��bX�t��fqZT��,I#b���T��j�����;��22u�.K�~|`��׶��� �#Z�����D������Yj�[$������R�x?��k!�_����5c�JV6�q��K�V�x[>��3��}����G8�����p�`ˁ!>t��L�`>�x��\C�T��A�X��$l�ª�D;���:p�Em5��6���F�_���6�0�V�����M�#�.L.��^��V�� R8�<���NgI���T6"ŀ0��()���g��b��l��qVoԊ��]<��X\ <@�A.k����Ojc�Q�����E��e�~�O.8N0,&�5K!{d�����t�օV	�l�+'���B��"u)�̏� :��K�����6��(	P��5U��3FP������� zm�P;�v8_z���8PD5� ��02B�R4�_ϥ*ST�7�6VXs_>��<�Lc������ҭ�%�Y��h�%C�96U]|3����?�4���7����{sW� r�)e:̹�?��.�?����V��c�Fn��x����32��F �P��`j�!I*y�t����}�.Z�cES�(1��+��ɹ�	�w�1A7�����ׂ�R�7���~�r���,�4*aF�1��J�M/�F�sk���t-w4p��yܶ"�;�LW��6I$����i4�������)��G$�_�e��[���!/pK�V�W/��Bܣ�(t�P�L[f^f�/�A�}�MK�TM���\qr3��j ����  ��
z�~��x���+�+;��@Vȏ[�UI9R�;Y@?K����p7�i[�*�h"�d��Ǖ�v�:):Ƀ�M��U��[��eHɸ�;l�4Jw�٬�	���@��KJ}������`83�m�y�^����&|�V?�&�o@C �\~��� ���MK�eD��[{N�MX��<��g�Lc�lG)}T]!_�x�-��}���L�S���8����E�Q|��X��F晵���3�EJ��K����K�r��K���x�4KX�/��Wk��f�EC���~E;Mεq�%��S�+<�ґ�P	�7�Ȃp�
DT�O���>�y��=!Rmz=l����s����Q���9�/�V���Ji��=�+�?�����M���im�J��۱�����`�����5;�bw�@��M@��BOt�fd�׹_�iW��$;�"K�)Qﵠ�*S�|\Bȶ�֪o��U+|&q�����ﱜ�7}��^���t�� @{�	�t�l�Ak���YfG�w�A��"#������� B�.�tk^>�$��?<Ί��?��}�K��izG�����C�h3��#���!�E%�f@ sp��˯J��1*tc�C��n�a�q����CB~2�;}p������	��葟��x����Y���4e;yْH��I��qN�U{)�A�|�]�W.��o��8���.ɴ�y"�DCi�5���7�`����he+��dAB�f��m3K%R�n/�o�~�/a2�W:��>e||��z�V<ԑ��s��5�r����u�'wE㋯��0�-�y������2jL�ܚi�j�{	ʸ����P�q(.����5q����O�t5$�h&d~��b�)�wVx@�k��`(������{)R��'�|��j\��)���~ə�5��O�(j�Ge�1�~�V�x�08M�.�Zk���-~[�E��q!t�#0�Ԣ>�B��ۮ禕��I^Y�ނ�k�K����U#ԣ�G���I����1�LTp�D%
M���k���s�3�u
��������IyM��p���,\���Y,�I�.�J
9�4ߒ��TҠu��+"in}�R!H��c���w�~�Chc�vYI����G��hŧ��,d��g��
��~���$�t��	�z2��B� :[�BO�,�ӞH[I �V��� U�ݹ��q-��|��Weݯ)S���������ڧSuy��brQP��/d` �T���a03j�3��J��::����Nх�0��ZD������R��9�iV`f\��B���P�����q�UW\8a�j��+��	�KtC q���)Z���i�Le��w��'�m(��Έj5���r^�Rͫ`f@� 㱼	�^b���"�$".��EMr�E�E�6�ww]5�J��~��-z�j�-��B�Y�?��uL�C��G�{�4x�0l�'��A��oP0&J��t�"����M��[0�K�b�(�M+qcH�n9�z��!C<P1����u�'���(P��;i��o+ER�sl���� *qVk��"EI�3+v`�4$J�Y��R�7���r���3�o_��u�]b&��b���({�o�,�WA���d�]簵0�R/	� ]�?�r����ȡ�I���w�`�`{������w��W�3�pK�D�}%R�\���3�3���,�◦�0�ȹ��Ĳ�C��Ϟ�'�y��ɪ���M�(p��Q��s�#�L���Mv�.aS��/ �w�' ��܊)��u�;���Rv��q�g��4͵����ثE?��Q�D���xe�v,��JKD��c�*��'b��5U���DN�sT}��&�b6�ɝWX�%�m�!��qkȲ��}2�bx#�X8�p!���p�O�$�؏A�q	؜&�����r0�'��N�&�e���s	;s��A0�J�~]D%Fi���9W�hA��/�-�X��q2��d�+�W���;5�M)��ɹ{W��!F�'+�H@vA������kd�C�BN�Q��y"��ĥ=�Ћ�+��|L�����m�E�_��`!^�O@���W�>12��b���i h���%B���b��i{i��&;���6���m�Ჺ��cӬ���p*���xr ������L����D�� Lʹf_�D����#񝢕cˉlƇg�~�]�l-�&���K_��)_��zڡP�ߚ��������� ����!`��jJ�m�@���~����y�/�HH/B"��9T�3ѾX��*�9S�}��k��d�+cLubi ��}RU�����>O��2s�V��)�����xBD�q�n��&���k��{�p��2(�����W�[��V�2�On�!�#V6� ����-�t��S˹o抣�rͺ���5��R�7��,��/���8��yeQ�'��+�ZE�o)���?�AQ�'q�wIp=1.�-������T�Ŷ�^~�i��vq�C�t��%{&�}�;�p}9<�}jW�I��x�wD������I�K	
+�AX:���H�XV1o�
���G0<��o߇\����<�����	\��H>�F��'F��>�"�0���}��� э�f�P^�E��Pt7@qh�<Sg�&�`?����3���?f���Vی1�C����t-|Sa�ߌI
�L9�u��D-�=2"�>_iؓ���,^
�č�)�K�7LG�Zp�]֨����{�v,���t��6d��+�=���f?����+$@����WX�$b%��-��E�\eG��H䰌L�c��tɍ)V�ߢ@�e:hr��-���?E��	�g�Vr#�u�Z�	2����_�{/�e����DgKG�wM�W�s�B�1Rg�8?-^��P���e"�7o������"��L��>�!,��!��~%O�Tf�qHW�⚻)��)�Ei����+�z���\�kKG4n^�K�����e-޺Ah���/X�{��o� ��#��}�v�𵕋c��Qr�&<-p����y#KЖ �܃xX�yP��b�xw.#:��9~u؅'-�z�
5��q��%Z�۠�*�I<����s'�+�dNp��7k��y�n��ݱ��`�:P��H�z_O��H��y�h�e���5��)�+B�G6�d �Ls^�,��!��ψ9xCz2�!%��c1Z4���r���@�_���k$	�v� �뎹�8r����{F�8������Eൌ����3��
Pބ�A����6�ĢY?c-{IDV,?,�w̶��}����p�"^�"��K��7�T�¯>��5�+�j*%��7T.�&g��)x��C:���J���{Q9���(�Ç�޹3��x��滪)k�I(�E�!�G$�Ak�M�nhd�H��b;Bx��VLb�6I�K�ߑ�$�
2y=IS��}�qz?�EY�:f@�VD��&9�8|��(�i�Smb0�X+]\���<��F �b׶�	�n.f1y�Y����p�H~,1Yk�_[V�J����9�(��r�J�����#�\�leƚ�~v��0�~���l�ׯ/��9:�HpE1��|�3 {\��_x�$SF>~�k)��	0��w����I	�/U �����J�xz��nw���W��!:Z�(������t>t{аH��?�������{���o6�E��8ԡ��DGl�k8"�Kz�=�B��k����n�n=IlPoh��	���V#g�� 5-��,�v�8'�b����H�|]�͗¿��m��#61��GZ0�95hG:Nef�½Rh׻֓��K�1�w(���s\�^��S�Äo0��������-!(w�鎄0=[��>�6�ǧȪC����7C wB)��,H��K��QcBAy��>u1�Y��9��k��*�HG�A\&��| �h{,�B�6��%�$��$����z����e۲�(>��ڥG|$��<�E�v-׮L�ؐD;�#�M�栤����4[�|�:�Y�ڴ�q�>�X��l(,���r��'VHK�ϧ��S~��\M��'�F�ٜ�,����P���+| �w����5^]�R��O��ގX3|�K�-���K�k����چ�I	���
77g\��ؖ_X��S0��.)�8&������i)�"��D�P�i���R0���m/�Y d�M�-���>ϣ��6y{����X�˿�
t�ݿX�(؆~��0.��!�Ж��������f-W�2)�Z\�OU���c�0����9�\)�(`j�<��]Cr�w��_��/e
䴻+��ݧy�R��u��q��)��9�p�e)N]��
���4{z��2tr��S?+<a<G}S�oH/!+c��K��Hܫ�E��R�Zi�os3u{F���閐(R�7���O��7?�[c�e$c�y�r��quI5j�6ґ�H-�L��5����@��BF� �zU\�:��`ݐ8̣�*[c����霷���X[�q���0�#PEnQ�k�����n9ý�w&�g%���{��֐ƹ&��+~���e��ƫo|��"�z�2E��Q|���ݓ�b:�K�2b�4�y�	i�9ݼb���Azդ�?�]��hRƃj3��ܻ&�o�uw�ç��bt U4�Jt�+�0S�p�IZ&��7k�i)�s�
[L%�o�aB�ϙ�:�}?����&�h���͕ƶN�C6����BI��f+M��]�Ӫ�J%Ep��s�_����L����{�˲�tu���cO=�Or�|�k/�`O)q&j��1F_a�����f~��&Eɤ,�ٿ���(�0���QL:��N!��N�����|���5v�p��2����{��r_���s��t�g��˃�(a�W���sc�t���x̱�k�U�`4&�z��}�׷�ه�H{�������f,��f�E�X�@�ZW�I�M�����)�3�� ��r5O��ˍ��P]˱J��$��"AO���!}�q9cı��J���j^3_���!�fӯP\�԰�p/_�f`�q�F���A�M|����
6��*m�J��u;	[�׳'�r-nsn3���wf��8U!��AK���_�K��>��?�m�i`�u,T)/n�?�E��^��&�@��ez40H.��<�Jwt���p2�h��}f��j݅V�4�YQ܊h+��yR�nm�Q�'&�6� rͿ:��u�(o*Ͳ��m^�{�X�K%��	_C�FAW�1<ZFvS3�C#02zM��s1�6�Z�p�q��w4*-MxDI���� E5�#M�.O�|
_�@`���#]v ��K���_�H�u\�_�>�!�h���M)�v��q �Pz�pk���z2�P"�Bs�<u�E�SDC��Jc	q�Y��I��EYj@���N�u1d����N��F6�c�|Uq��x`i*q�}�,����]&s�?���/y��Ysb�� �J�R�8�s��M<	m�V�#�S�����t8\�*��kG�xl�k�b����WH�)�ןN���h�&���G.�փH����7L�ۖ,�~][2m5���Q�-	Dl ��E��Ư�F���V#����z<��yMs�y�N#����;�+@Z�R�.˟^`�5�d��4�����2��������AN��c���)��z�F����{:vP�t��@Oژ�����=�j��Pz4���� )�X�K�z�X.w�tޛ���O�v�c~+y2�����I���&N�?et�գ�e,��&�p�X��AVߌ���xTF@�k>�П�5�ь�t�c���Fk&x�m�u�����j�zz�^���rЕ�BH�#�Z�"�q��=�AQ�������n�O"�2��9uo��]�ZV��Z��M�H-^��C�C|B�	�µG�Zӻ�u���E��K�@&�G�Zˤ���q�=k��(�g#c�I7�R\�K�.���f����bͪ���m<�:W} ���f���ް��b�*Y��Rc��p�q�B��ag68��J����w:�vEx��iԦKl}j��* i���1��3���M�hh��)�)FW��VΞ������N���ɐ�8���=�#ō�F�U0�/q�@u������Pv��+�/�w�Ѳ��X��ۨ$�F��\o~Q��+�B��`�x�q5�Q#���iɶ����1��҄lp4��W�y��r9�t���yɏ�Ə´��peB�H����k�9�q�6:Gm�:	�ޘ�W�����o�(�|��Z��ä����Њ���v�XH�Z�,l��d��̫�^�4#%�~Ab)+�]�Pl�$� ��[�]��Z�+�f����Q��U�������q.�oA�7��:6}�CCۯ�f�M��2q&�O�  �����@�����g��I�ٕVs��n�-�>׊n56�Ş������]�$[Ӈ�*�����D��I�x6ȳ��UB�3R�ϙ�TM����#�-��v0NI
�;�� �a� �������"7J����FA��z�#�B`��1&���q?�*OÑ�x�z���g,N~�ڕ'�H�S�hȣetكG�gM/|�r�c�:�^h+��T�J�u�H�4�
Y?��/�H�:��|qK�e��L �+s�rM8k�V�9��ko�2�q���.���Zsv֝!��:����[խ�^)�+��84���MNz8It Yt�^g-k�5�4��5���ޛ���2;�j&��i��\�r�_���fQjp�
��Y)�f�-Y0�~qr�a��ƽt�+��-�c{\3��2�2TʛE����6�pS���̮�,r	W|��͝�7�q�,�ŠP�e��y��=g�m�N���T� E���.��g�Yʚl"���3ꮩ>���$��
��c�Wk��h�I:�U]�z1S���(U�2\�"^�3& �+��p`g	fe�Lv�n�ۗ7��.sse���r���6y����6bâs�n��|!�scKh��i�i��v��&T�dΑO��Ʈ�,	�W��-,mBR�Á�>Z���#GJ� <]mcXky��5�^�qCb�n/(�s�P0��Fл��x��B�q|K2:-�ᔺJ:+6��e<��(�c9�5�J{����	�-�68��H2	?���e��Z? ��7��n�BE�g�(�>i#%�P�i�3$���c{ݘ���f�*3�YJ�\��o3�w���e!�	e��G��)� !�ۛ�v�~�0�����M'�E�|���c9͏�2j��j89/4>�v�.o�Z��1�ϐ׃��KZ����X���iE�l9�����s�A���$��f8�t����Rq��M���^�Y/ʛ���1]��V
��Ey��M���vŬ ?�c�Ȣ	d�&�.AƐ~��:(Ξ1X���_]�3��������'�ˁ�Ռu��2�HHўU��U�s�d$ht�yb+�b��+��W��3v��n��� uaoeC⮑xe�ܙ#}A�ma��SXD�o�0$�_�)Q�(���0j���B�4�d��޷�K� �֭�ѻ���M_�����$�m5l�eO9 {�1�]�:���U��YD58�Pu�"f~nn
���ǖM��;��$R8���9v̩Xh���r�=k?uШ�vpD���M*�&A����"5JZ�6u ,zr0̈́_ө�m�n�yP� '����
eo��#h-�	w�ːI]j4�e>���)>�k,��#�ܬR9.������nLyK/���Kh����r��3ۋ(�%���S�]�cn� NhqIN�C&��*굶����lU����H?���z��k�%�+·F� ��x���Ur3q��Q?�I�z<���V�|���o�Wl������ �  ���s|KE�(�4c�~ɫ�g����b%��V��U9u��1�y����2���	=>"��%N��6iS�Y��@,,�N�πd�����l���g*�`��-A���j�e}Y�jqДǋu����:���=��ǘi����~ Q�� V����<�<�~���j+����cTϚ�-��u�:9�L/��#�%\�&���u'��]>eF�6�4|-����D�RBF���.��>%�����e��tvb�6���kǻ�I$$8�����K��?DI�EWăH.�)�ʨ�6���Xu�_��g�7e��}�cI�0i�<o�Z��u�JҏAkx;yٓ�Szm6�ct��MD+�
����>�i�m|f�#�AP��39������sR(��6�u��T_��A�͢$}�nXw�(�F$�ʯ�f2��啌A
�MФ�@>��#�~LP��u1��G!9�Nx�I��&}�-��;J���>c�<O�J����ɝ�!x��	�R3Ԥ�$����������&c��¢�;�;�[�,[�H27��~�Ŷ�+�**b��N5��1��hvTevO	T�B~�ڹ��}M��)�l��Zf_��"?#P_����V�9!�y� �#�y^"�f �,�b�}EI߯$��[F5V� ���3o'�$\|��:����F�d�������bk��)�Ol(7l��i'�Eٯ���������b۷<����)��b�" �u�Bq��M������W��Ͽ��; �nRyYp��02#�<��/r��ә�����F���g�y�B;�?[�li^˷1L�$���x:u4��mŦ6�$7���-�A�g����KR�DV����U%��b��b�������kd�?��˸	/a���0$��h`�Ң��w��T���},;��`�=�h�u�=�с��,x�Y���7@�L}m�ĦU�~M7��YB$v��`X��Q�6#B&�AZl�h(����E�窱�Ws�	&oXf!?3�|V=O7�,�|������j���@�{����$+<h���x�� sl��	
)�VH��F���F��q�����Y^-ʍ�NX@+K�)��⾭�-Q�fE�yi� W�I>��4t����8	���-�{����̅��`��#{H��4����U83ˤɵZ����H�	A���m�সؿס־XX����]�����)����7)+F���"��C��)c8Q� �W��z�&p��f*j����O[{����t�"u�f@��7Ul��:�u����앀S=���� �;~�!�tD\ 4��^�y��H�fbk� �z��6�$����C�v8c�ϿT���jJi% �n�]K(�qi���d�3Ϩi�U��/lSPr��H�Y/}Qۑ*4!'G���JWF���M�,�*��㎟�?{���uPw�AML�����hFI��a�Y�}��3�b��F���D c�\��ɟ�Ű1�� ӓ����4�� �� �+U�s�N�?>�|�ƚ�=NEA6�9�4"3X�)�'���菭�1��J�{Gj5�G�HQ2P�`���Z�������p�攢���\�8��{Wr�:�iZd�9��ջc�O�;ꕈ!�Jl�aCH��ނ���ǋ,q~)(�8VQ�	�	s������˞�ʧ�A�L���s�弧l��R��m�C�6q��4���,'��g�%�M�ZC�� }}��]���Ƥ�1fU��� wj�Q�Wu�C�1�~��ڍ�>��;zaM�F�y$���\y��^���.���q+�J�%��� 㓑��\�#k)u1R�+^M���/��-Q�t?�DH)��֏Vb��,�x������#0��*]^\>��5I�Ohw��z^�U
�-Yl6�*	�{�8��h&����kM����[�Ȼ͊��*[ěvT�Mz����7
�)�aw��g�!�ǝ�fX���N=Z��/��j��&���߿[Ȟ�y�3wxo��e���-;�Ơv�_�A�v���:Fi��U��%_>�L�_G��&&�`Rm��Gs��}>�kGI��J�&��_�	�f�� ��G?������JU���X����z�"Q�"[T2��_QpH��ֿ�?�3N�c
b�3�EBzA�;�mR9�;I�7Y���?���$����\#��,լ(Ý>��Kq�uOz�3E$�o�ʊz3�B���4HCl1��A{�\����z��d{ŧ��Q�G/�?����#�Dr圃+�iIU��E�0���ӓ�k��"�%�ʛXLb�`�$�JK�+�#�W:����+N�,�����C'�KP"��S��@��Xg6�Rz�se?��m��s�Z
B�eG�辴��N
b���j"���k)}Z��@zVAK5�y��������j�xư�����1?&�X�'˝5����|�\F�@̝\K�	�Hv�o(����cC�hL~K�-��C=�P�c�f$��`A��ҋ���B���V`�?��)����$qAOj�$�<�k����5�oe;�9yß����D=�)2�]�~Q��a��S�ņ2��ط�}0b�)�GU#AR�����.w*�G.7�s�z��L#��&�I���wh�3p��I㗓ǫWZB�>$9��nđ�!-���딊���S[=��	_]���X.������,�����-��1w�,u`�&_+b�����ٓ��bJ�2��y�1�E�sX�S��<s6̒jk������YA@
��F\��5
��J�×L�P�2�_�&��B�i{'AD'7�ӈs��ᘆ��RB\bIO�h^�:Eլ�\z����X��^��h�F�[���]/��,�W"��i��诪��
>��:Z�S�o�SJ��i�����|]�(1"������U�jw2M7{jivc�|�;�+��I����Y�Lyo�b�[���۵�n���;=�ۼm�k��["6�D���/}�T�l,LU�B�(h���/.@©�8�H�u�evuL�0�B�����d��G2	��`wXU0���@��'��O��ɀ"�l5ލ|��h+���Wߜ�����ϡ�'5L�͕��`�L���cwc���>��Tif#L�y}/�9ݿ�e����������a�i�T��̤n�6�E �#�A�
)��=���9����	��&���$��U�=A�B�Ϝ��j�},`�x�Y> *i�,ҭ�v�}_y����qNw�x9��<�R��'.����|K���s�+^��n��bqIsƷ~�?>���MZ9������֢ï竪焍�!c�v	4���~hu>�*�wu� �Tk�|�I�ba�0w>kI��.���^ӰkkU��wU�j���v
\�5)EY4��P�w>}�$d����43H˳�|� �Q˧{�8���n�?k�L�&n�7^���7��4������>���//B@�M���L!���C�4J�rO�6Q´�n7b;!$�s���©΢WuR&сc���τh�B����J���Ð ��������р��/=�YH-C�x�N�kYG��gxx"�pi��˅��o����\~�� �@c�N8�",,�)�zURӦ:d�>x�]�"#����!�G������%��zQPÊw�^�N�cg\Iˎk�ۍ��v��# ��c���h��L�a߱���HXn�ULyh��5i�ɝ�2Wu[����ulJh66��<�L�R�%m�Z�Q�G��Lh��=\%��2���tn�e�wN�>+��E��%��'�!�K�	�=`r����蜯n����<�пP�%�n?�[�����e�����R�+y��ӌB&h���|����yK�:��|���0ޓ�Q'&�o�n��������u5S"n0��꒙I��i�e�M�H���������ئ/�A�9U����U�4[�=Ud�Z�&��7��ZW�{_i��/70C��z	���~v�Ջݲd��QAv+�zij�V�z��Uj��peMtV�z�ͪO�@�����X�54�=|�dz�:��_N����h?.-����!.T�Deز�8OHѽl��,b}f<z}�:̦�X�Toi�B��ő]/ ���G�6�V?��l����uC�Wr��r�u��[�e&�F�Z�,H���o�m��\i]ݶ�ZYS������7�����ɶV�I==��o���۟�S�����_Jq���lm�"t�1$9���j��/��S��ϣ��<@�7 ���}I�۵X�B>h���5��?5��&fO�6HLx��6Q�8����3��>��d#��S�� K�cr������m�_�[M��
�"��oXH]��B�qθ�ܶV��N8�Zן��o�����R�ҋ9�7�#hlZQ۩=�Bbz4}�z6�>�TJ1bi<0�[{���w�WZ�l$�\A�}�~��>��͆�R�,n2��{���@v�� �D*��Aܸ�q�K=��O]S�x)����MM���q��m81��2w��z�&2,�d�¿��@$I�a���z��M�d�K���&�<�-+���(����\��}��qH
��F=�D)M?G_�颏%�Z�Y�Mw�?�v6�]���j�	l\;N�K�J�L�I*9y�b��F��1*�)��\Q�F)e�cmN��<�i������p�L�ܟ��{"��8�����vr%' ���ß[!,pzNl�\�T��!e�v?J{،�(J�x�b_p&���Rͭ�^�j,>]D2�Z-�Y al�9�$��!,

Ų �ӷm2�O�q�X��YM?S��C:�zbF���i{�w�n
7g Z0� � ��v��y~���ة��i1���o�V+gKѥ��-t�y�bxU���P���:';�*�m�N��/->�{��)��[�����T�*e!3c:c��?�͐X��5!:r�τ�d%(�����_01o[���B�i�&(�-��}$����K�2�����4$Z�������\��bo\6|�=G���=��)��I��|�V�8\n+\4�OXO��m ^��[�#s����&�p�)W�{�㄄+~�n/�)�Tˠ��a(��,P.0O�k�ߏ���gTy����dG+`��=d�����/�����)"��,�a�����k�@+t0�@?�+����*|�E}\��xh��M�����o]�����)c�?�4TI��/�)����n	5�@��x�׭���(a_�a�Y���8� �"�]���J~}�Q�d�VQ1cOT��˛�N�6��C�0`��9��lA�Z��hR��w�K8������e�;��6��ޚǼɰ��W�^�2���#t����v��
�U��f<�/Zw7�@&�eI}Y�$�o�Ğ�|c?S᫤sP@Evp�%Ơ��^}��>ha$��qТ�I�^9���[��?sҵ��֎I�����#��"�X�Yk@H k
�m��Q���V0DR�@?%����7��> k݉7���z٣����{A�o8v;S��&I���c�	Tj���+��r�x��0���.���:՗�>��s�(
��O�xK�����d��[�Bdt����Ē�an � Pz���<�
|{E`�iSF��Š��>��~L5��U2��O��)XDYq�тoǋ�ӁCJ+J�AT{0i�CTȧ�I�e��?�B�'����It�X�@,1���U����#)U�n`�"-�,�%���v)vʽ�.K2�����5g��á�Ŭ���:��/��͈[@0A$�I�-��h�rT���lX�P�X����b�-�����G� �i��j���^U�W�~�[ˏz(��C-.Ky�)���ꐔ[�E���7.��ק�+=��l_�_��I�vG:ӯ����b<;ƪ,ˁ��_�f�zbD�g��ў<�E�M9/��$~a��\24��k��0����Ձ�QW�yͧ���gޝ��.�rKb	�Z!_��oj�8�������I-?��"�m�ѧ���d<aQϺ떳i���[`l�i�Fv+,ч�b{p��_���7'J����Ĭ���%آ��Œ�BC�E�h��٦Q�	I;�W0~ 0�E�� �+w3���M��hnf�6�hPy�o���$�IE��f|������6�����^Y�P���ߒ�ώ��NI<�;\uCEv/��{�P-��R3T��i���8�@�)X�����4�S�+ۅ�;Ϟ�_�W��:�ݷ�j�����5P�1Ť,L�?b�ز���*�r�Н~�Dh�6ݰ>��R�?@=d�8i���(�����"�s�~w���>ث��*w��y����'��޿"�j2�=k�Gzb�����($`Z��/�-��Rc�ٸz��mj^X[ʎ�˽*W�N�P�Nl���4�&,3莚w�:�%k/�|kh��3�XUe�����A\ʕ��B���:�[j�
�8����� �ՎTTO���l�O�:3D0�D
T��3�kC�ۍ���VXq�6s"lY�,p��d´HW�D�����E3\����G�ք���<b'��zκ�h?7�����-�^��`=����V�à�5��'�Rp4�n_�[q}���G^�d�����ȃ��2i|E�v���<W��^����lYk0��\>��/�9�`�zO�j/i��6]k��j��4�����Z��bQ�3Q�%=Ǔ+o�.��"�$�c)��G��u[!�9r�k7]�Zo��)�aT�0�Tu�3ԍ�_:B�m4�I��e��!_zf�#DrU����g���t�W֜���������b������aE';� ��U	���L���sO���gOkZ+-m�bA�f��nd�ő!U�cvH�5�����V$��`F�.kQU�
��;`4�i
O?�6t�0�w����4�����J��ɸ�p�
7��R�w���	e&�!��2#򯱐g�tw&*�,װ#����>h�ŧ�~�gQ�{Q� �.;��v�a�l.�ա�F���^+��C���Mi�Bc�7��(�]�cSky�=��fǸ���m��;x|s��)U��Wțb3��y�ߖ;ߪ[�R���&�X*���gh��΁�7r<���
D�ѯ��R�����d��F�A� ��U���7J�&�9��6̀����,��E�O%�A��	^�5��&k2\LT�N[v���;���-�QJi!ĺ%���"�f��`��� %4h!�8k�0'�gkϒ�V�o�/������6��j���W�L�]�=��	�6���}ʩ������lj��(�*Ό.E��^8�>{O�,y�	u���gX�2����=z��	ΐ�a��!2�%�Ngn��C�z��]i����V�?�s���p�:2&�6Y"���hm�o��K����p˦FQ���p��tt`�#�%Z��s���YL��J��Q�[�}Z|��r�Hi�BW�$a4���,BAr(Z����5OW�@��D	+�v
�&���x܆�b�+��b]M�I�r��IsgkV.�[�y�0�a���O�;�Z.�t�߃�W�����l2��^�*%k��� �R��qvY��YC=�$:(�b����M1<$�����#ȑ�f.�(���n�gm+�r!�^;�U�RZ�7��$���3O�A��c�6Q~v<���QgR;��v��m@�ɕ�h�~��3����[����4@V�38dF<���BN婆��!�I3ʊ�=��~N8��l�	�s����oj��Ep)FP�=꘰��Q%�7��URi��~�Q1}���7���ޖO@D+I��m �BpzL����M*u��Z�3��8�&�!���O��O��T� �b��_����q�����zEL�D��1,���#��kyI��}���O��i�6vh�:�"�K�>�b�b��I�Īh78��&��	b�L�M\��'� ��0��_=�=�t��}-���iz_��_��}x0ُ�C���1m��}��H�����I��8�{�6�6E<�w%L�f���=�u��O�,Z��O�uba��t��I��޺ME����t+Y:�M-��.b7�C����j2Ch��F����YZs���W�Z#w�4FD~_Dm���;�%�L!_���d�Q��d�~�q�o��܋��Bn�ڀN�0M#�0ߟ*:�'�ז)�u��t�K�z�yUE�oi��8@�1�6�N5_�"��vDO�m�4�t�&\�[8��#�7��L��}�zP�*�1l����������(W���-��<JEpr�0����]�G�lX��ubm��oS�F(��~��̗=u}ͲXFb�E%"��ֹ�r�B��xs
E�����+���`)+���1�E:5�M5l�8��4��WB:�F1c�$o����s�R�m9�0!ҤV�B�yV%h���6Yc����!,{��3]ýd��$�Xe�N���R�<��P{q���1Q����_U	�j5u+/9!22[m�����Ҝ%���i"���3�9��c���=F���غf��@�lPmU��%����8g��V��/l�xGV��k)����b��ֆ4&R�z�4yf�~t=��$��#��z�AP��|�^�u'F�8o�=/��S���`�����.�x(�$�N���Sd6����S��-�p�{�љWD�a��Sa��Y`���w���#�^�^�D�"@o��-y-p��9���>'_�W���OݳX,x.��?�}
�1B��%�l�aw$[�������2ͥ�T���Y�w�TQ05{����Pqe� �T�v�� '�cٱ3���?�JJ������@�q��W?݅�����y Z��x�t���-���'���@X�����ʁ/������
uQƫ�2E�c�y���iB�v�B� llfAg�Ig��cE_���I���1\�H������`Oo?3��U��UF���,?K_�iW�Vy�((���NL�?����y3R��ϜF��N:b�����(�e�S'ڼ�#����q��2$N5M
�i]rd��&������n���������KvD��txv8�*pV�hԻ��x�>����ѝ�!(��sq5r;�
�\��C���tjj���!�l"{���-�~�lg���|��l��!B���<��_�j���R�4��(6n݀��yBV&>�������o�2n�������2�2�Jͬ]o?��J�AH~5Rg�Zh'��ZsU\{I�����q����]L����g�5b���f�����FO߫���-��+�Z�;xw[�,��c�7`�#"pЊ�I�b*�x�>I�u��c�|�k2�Rը�
� 'o��\��W���LrTD����-��+!d�D�K��0�.|�H��s���>���%ی�|W�@C; �y�Fi�S�o�Ю�,�����K��*&��;�B)��	����� �u"&�8Ќ-��q�*���E��
��ni��ɻk�ΣfU.�/F�Ѻ[U9;.�X�6ԗ*6��Ϧ�a�3��G�8jY�׎��U1E�i�2�����$�$X[!q��%Y��x���-�0E7�f�7�`vhx�4���]-P:~[3	s����!Fw0{������u�1L��@B���h��� ���|�d�H��#wlnG���J�Y�$0_22�ə6m���Ĩq�	3%� R�{�:��b�r9��D�e]�X�=y��9" A���-U'o�¤㒭${6[��.É�L�����h���Y�x�B���j�r2�1�W�w�L�S&�����ͨ���t�� �.
XlgIbX*�a��3����|Q�6&����'��T&��T�q-���h�`<4 ]�؈ޤ.����G-��5���i2y)$�s�<p�^j�o�������g�޾zهBMt�RS�4[/0�U��P�W�M�����@nC�J��RfRj�>|o?��T����֥n��H��LEf�+�H� �JY#eT��j\�d�`��WU��ǲ��ɍ�%Nb%��$�)H�	�GtJ�:�5���w����;64�	/.
��or���]��U5 _LƞWԫ.<K����9�z���ܸH�	ج�gO�5��޲|�K�b�V�߶Ɖ��B�(獙YR(ٱ�����\��ֱ���jA�D� �Xܙb���.$ w*>⢶�:��g�Bd0�E��B��S>S��Ag���!��OGp�v�a �hdQ��]�N.%B�f.ym�~@\��%�����x��8j��M�Aa[o�e��$8n����v�g���0+ N��g�~��,Z8N���Z���0q����(ި?�(���]�+b?�n�����|�#��nfd�B�E&Kw��TM�p��Y��d���*�N Ŗ���,���Sj�p,�#8�:��u�_�.������a�<�$[ų�ߡ�)[9�) ���c�r� f6�4#2/&��)�&i��\'��Q!�y8�| ��>�n��i���x�i"��ܹ i�-
�{t�~ʹ�ֲ�u-P��K7Un��SrKZ�����FP���@��]�%'��{L������C�!�>�!�0\!yD<XZ�%��ݼ$��6�'!H�u$�Q���Wu�=m�wY\lh?���ُ�lB/*�o�bv��S�w�5,q�l
O�H��l�z��5���v��h�l�*�CJ>�
��'�c��'�J����n����B�.?H�����4c|��!��^,�����	!�������ǡ��̄M�9�h��jm�1��1c�8DC�E��A�*BС���aǗA�!�H�@��$lrA`��`��̶�3qM�k��f[�\Hwe�M�!O>־o@����y�I"������9�0������'�8����~��c��r�����k�K�@Ci��^�\�������FD�>(�{�5���3�(�)�d��&��G��A^���FJ�+h%��WV�*.s^%��ac%�	!�7{��UhϭO��ey_��m���W+�K�+�YEC�� F�^vnx�ۧXU��1�s�.��3F%%C�,U���3���,j��-���a>��d�����5�h�CZ��~<�{ ��L답@b%I���BB�Sd"O�xG��n�S�J���^�P��#���Ft�`]�}�n�2���sK���MQ|(F��T$W&A�T7�_����ݰ�:����w|�~D��\M�W�%�Ө��c�����)�;�)���imxτ�Si,=ݸ�kT�>m���~��b�t���3f���B�>65��N�(�k٤�)��`9a���&ۙaq匛�K[����ݖ)�a԰cn%����џ(
�cD��5A9�ş\܇Q#<؜	wK{������t}� �E|/	G3��j{�9���y�;{
�B����s��L6�9H����rri�,�B�a�ݿ���U�7�|�������u_�A0�N
^�!2��1b,ow"4��&�m0�|UՍh[�j���]�UK�eY$r�}0��u0j�A��{�sc���<["�����v=0������C�X��/CR�%Y�=-z�ޘꌨ��nUo�L���sY����P٬��
a�~����a!p�q�ΛOh�^���U+��%�.�m���{�^�/��-C��p"ТbR^WZ�[����قe�k������T	��R�5#_���<oJ �C��(�@fI���}?�ZW���ր���:����P ���΂f��p��,w?��n�(uMz�����!��{�pA���.�BVzC�>C0j���o\S�l���m��ܬs���1#�.��cɨ��|��bOe|^WyT�@�7���UC�?���p��vm�c_.3�o�s�~�ʈ"�^�l�+Ez�w�L>w�	\�*K�0���A;�ߦ�8H���O�%��_�by)���X!���c'�~L�̇����h�	���3����U/�D/m;L>1D3����;O��ܿd ��x	��:Ԟb��&�a�Е�Z�UăP8O�� N�2p��y_�����d/�[�G��I�	&�Q�RsM��5y�@����tt��Px��̻@t��EV��1��3�Y7�EƇw���4.��M2 QD�K�^ɚ>�*��0��Yͣ�QQ{VN%��F�@���J{����������ҟ��q������F���N��sm�ˈL�?�bx�p�sbOڲnsl����E ���C�!�T�����"�3Y;%*L.}�$����l��ѵ�QMH �AGv�D"�կ<������'Q�iR��|� c�(,��s(�ؿИh���$�0�aT��޾0�	Oc޿��\��F�d1 ^XT[�	٠�O�����_S�홑��{�V�`wۻG�����elvˑ]�iMRrxZ��D��8�KZ/��q�X='@��`% o�e[��]����4Q���ktp�A
�:O���]��\��,�#��N�e�G���=��JIT�DA��5�Suv
�g����O��f�+��tB�{M빁�M<�dF���L��]h��5'4��S$F=/�E��(��Xw���f�<R#�QK�YV`��:z�a$ ��� Q���R�0[��������	�Uf��o�g�2=pN
״��^H����m�R�>���R��v#��I.dK���Ď���@D,��/g�0/>�i<�F�v�ꇆ]���'�b��V�g4K��l�����;�9U��
/��s6�APHi�p��uJ�_/�ڽ��h��W�t��K���۱.�Ż�.�yRY>E��@+���,�B3,h�"����$�:kq��D�+�M+�򸗛��>���$ ��@ZeY��v���<^,��tS�%ATz��|�����h�B�4f�eCM����e��^
���Q9O9��&L�X��.�4ڴZ�r1Y�%�S���A����DiZP9`K��k*֤�e��E���?� ��)W��'��`�v�U��Xr4
�	ۙ��
6.HLT�#����4F�͒��+��`B�����i�d�g6�.+� �C�~�C*�d�s�qUo9ޱk�I��)?���Mɚ����NDYa����?B���0wX�c��$f���9�Vͱi(ÝN�!Yv�D1� *4��v#�~z�j��M
��C@&ٽ��;
i��M�ڨ/ApY�Zw�h�)���s\t[ �)i+n�&6��P�[<�_o�q�F�ή:И\�ˢ�^�z�ģ&�UjxB���`�1�\h�����[��>�T����=��'~o�6��Ia9'�?�A��vDqx@=����z�>Nf�Bq|K|c9�;>B����q�=p��R;-��u�h:������}z�[o�-J������Z�����E��;,���^��v�R0��8�[�ză��ՄX~w��N ��;���(��C{hP?��I&�4<E�f�ԫ���6b���,]�-'!]�����\nY���*��}àrsx���.�I�A33P�Xt��O�՗+Փ���;w}�FG����]N]a�G���m�|��Z�a���HRj���(�	�J���iH��A���^B��R�_*^��'�`�:ȵSu4��}���<#(�ˮaS��/l��r8�%Z��#��Q��	�F�T$1dKr^K����P��S�oE|n�V7O5_K��w�Ɨ�!�p�1|������5��P@��i�;�����؎[c�q-�iO�)b�p{c��:mQF���C0OA�g�
��y�Z=d�_K���}����"��,��0���C�U8/>bp���ƩޠU��C��wp��M�-tw�St�ڡ�~N}zK�HP�w|�f����U�ةT��D�aA*�� ��,�������׬Np��n�4�٪i�0׼�cm��֮���!�/�?���e��E� ^��Zzw�Xe#�ـ1����[�_��,�3�c֤TU)�7
6��X�V�\Q����<ե�i8�6`����v<͈uB��y3w��\Ye8e�J"i�&$�[��]���保�Z��8�d%ss�H�9�O�;����u*S�~�b�.v����ӵ��5��Y`���F��ZdQ�}|}�wl�oڒ����m�Ubw�\�vt��	ނ�)U����iu�h�So���Tdq�0Iw2 .��α�I��)�g������Lqv��ٌ}S���ǣ z�G�W����zK@R���_���5�p{�4���ͷd�$�<�B��*C��ii�*S�0BC�-P��|}�쟥�i�y
�^�o3�5��8�#i���|�$����V�(�5��
��p�%���e�S����/�JJ�=��gy���h�Ñ�鍯(p�SJ�N.��&���U��(X�Y�
D5��ܿx���ed�7V���*�RE�D���Y�T��[��h��]���4�b�:�- �-��`��x���ЗhؙUH?�V��
CT��)�;�*8��Y�5wĠ��N��C�"`�j�5�%��C�<E^�NvPHN~����� J6����-�>��/q�BQ,�瑓������N�TӺ]�m�U���|6ӛ��2c��B�����i�ńE���yP�8anS)�lp*���s�M�5�)��F�f'aY'(��*I��Cװ��h�a�pG'"�`p;��"C�;~+��$�E23�"��*+�)�I^vTwx�|��k@9�y�_YICR:�/j�7w��������^��2���%I�ZdᯇJU���F�/�C��t�)��_�S\�wT�ej���ԫ$�nw~��JP��C8[�/�^��Xř}�`O#��ʩ��vz ��ŝ�u�d����BBٲq9�@�K.:�i�J\��h�Z0��]��DˆTq�RMF�
֠s<��K���¦}�i�I����zۂ	�eF5�@H�&t�&�-J)�Y�_NG� �j�Rk7{��!�iYSb ���i��pҲPI��!�1hn��3�3��B��D�W��ZxC�a�ຼ�¯����z�[a��<��ֻ����I�r���85�ъ�D��I�� �����n߾,kH�aDՃ�VУh��=�. �(wX�������p3=��X�� �Z���D�G�3����L��#�%��M6Ozj��9@ۂL����fq��ٸ�v*�#Ũ�` 2_�f���ܦ�>�[Tl)��u�E�������ǔ���`6o(���O��/�qlLI1��;�Ɍ#x�Bt��Xai�FDm�HJ��c�S����YJ��6���1�����<)��/���@U���W��9>W@��L������ܼҒ-��>N
:��ASC�)wf�j��#M���Q�/�I�=1O_�#��<���t�5*����7t�t)�
\i#a3��	���s�N�Nίb�EU]X�	;%�.�׬$�k1�m׀C[EA��g6w���L(�h$�΋�@6�0=��߿�F�P�(��ɖ?�d\��EֺL.��}8�oa���URA��{�W����g��޿{�hc懋m��WW.v�;�=�u�|C�;��=�8��\��g�t
�/vK_K{۴�W{�5��63�~*��h��������R��a�efgk���#2�z���������4<����A��<�;��"��W�p��` 5����I��<����_C1����[�Ѿ,\�B��{���&��JGM�opxR#7Ǘ��f?�^k�\�=�O���MW�ѣ�x��p;k[`�*D�meY;�;�ٱfY�N��5)�b�~��������:� �y���Ճ�\ă�X������<��. Q�i��6hEƱqe�ƺ�#�>8��%h�]�
o~@�:J�����,���@E�2s����Vk5#\��쀅T�V(C���}Co�6�^�8Τ���ב��>����<l����񋺀<����(���S	ܪ���k�~�8.���˿�Ȏ����ȴR�{����S�g��)��7�zjrI�s�+���
u*w�k������ێ��H�j�_����ι�}b��M�����
�D������wL.��b�qU�K� J�c�C#�|ӸCy��K{�T^\���0mVI9ب���q<Aq�]zOs3�Wȑ��-�s:K�����#��L�� "n���t�b�7���@c�ݛ���G��+~D�qrGMula]�Pp��;vگ�����Ş�q�k̽f'·E�&�n��j����"Y3(a�eSU[��V׫z�9*h��˙�ɞV$�Q��`�di�%nk�+w	�2gK,�#/^�*�DLH�S�9<#e�D�	�UW ��٭�!�ܖ�w���B{R.WcjZtN����T���D�,O�A� ��`��~>�b/Q˲��|+�x��9�Ol8ٜ���>R_o[_���i�v?%�z/�߻<g*���k���&���~�����k��Ï{S���2��e�|4�!��yǴۍ^RM'��<�[X�n�����.�Żk\t�QEj���CJcv�U׈�i���af.�^3�����U��{��ܿ�z,�H^�F��D�,��?����]m�˪dZM%��qd�Hs�{��K�m�`l+�PU0�b��c��U[f<�Y�N7���%|�0��G���/kP���;��tVŕT�k�����8����%Zg��Qp�uș^�Oy"���f�53��$�8��O0�����(������T�)�;�8��s
I�CT�:�(��/w��>Κ�����|����U,[p��kL�S� ��ێ�oR�LD,z�S3��}_�W�̷�+<W����-)�@Y���JӴg���V����nӬv�}Je/ކǔ���g_�P�{� Yk��k��C
/)�\�q-��<
�C����'��W��qH�!�W�q�� �G�U���=������`X]�n&�T)f8����G�2{S�`���Q�b��ME��>B�*������(f>a_�
�QO�v�����u.(FnᾹ�0	k@�b/͑1�P%os�P�X^v[��� ,θw'�8�)�I��v߹��$à�a�/��1\^�A�eh��?|�Ŗ`�[�[o�V�Kp������ɜ*����w��V��L�@5^#�T�Չ�{�l���S�Iiꛉ^.x&y�5I��'�7�I�Ck��~��Pchp2��q [��ֿ�n�1z3&6���i!�T��E���|�;�S�y755h9��	l�C�!��rX�^=�c���X�RO���U{��?3�6#�ɫ�T�&�]s��8�H[pt�fC�\7�/<�E��
�K�1i��K"�~�1­A>�#m1{���eD{�6#�2���m9,i���I��d�GMw�_�p��RD��W��ʎY�p�=����q�ON�r�8���x.��H�=��P�����|f�r�fhd=q�����+m'��g�\.��ͮ�;�_����J���a���F$�J�!#�o�_�kq.�i�0z3A�b�����:$�j�>��PEX�'N��/6z#K	@�+hl��������5�Qr�����^?n�͟H==��p{��K�M�=�"e4*��kyV�����}	e�q���k�O2UMQa� ����e�RX,6ڤ�u�g�����ܞUq~��
�����.�Qd���hl�p9cB蒢m�jE���	 f*V��ǵ�Ffõ9fe�m�
���;�0�
��wg\�$1�D�nn�p�p�x�ڥ�����o���m;��ku{j�xL���1�����]����Җe������-4�+�>���2ӫ�W]]���S��>�)P,|��<	N���w���w+hi0��G�)l���?��&�˓|t�D��x�<����0%0m�K��?b; �˼���jkxNS9��,�r��`p��%YB�a�!z�N���d�"l5��=��;M�u+��#g%ӈ�t��Ϝ]01��<0
�Xn�)MgG��b��� �:��f˶u��j��Jdѐ|{�8}R�`�F:�ԃm�����W�w�/�3f��/h,�d��|E�r;���M&�v��rJkA�fcS�!�D��d�l�񣐪C@�j(�k�S������+��0zAT����n�c ��T D�&۫��S Z٩}ļ�HS���Q������r��f�]/s�-�6���R5 7EPw�D�2���"吔E�3�mkT=U~�����Pw}�yj�:r��e�!�_M�S�T�~�#eNh���I�h."P��h��İج%�<w&�+�-���ˉ뤩�,��f��u�Vi]�	80�+�Jڶ�.L��1JM_�5a�7E	l�������DI�9�Y�\[�.���_�8-(0�\��<!��c����Z��)�p�i�+���o�=8�d_`'�)�������lJ�����}Ҕt	���⧰ć/�v8�g,+a�_g��9k���[�[�G�z�V�-�Y��&5�����Χ���h�.�y��E��U]jg.O��(a�bj�,^�_OVL�o�Hc��O�0S5V�b۷G[��y�Nj�^���se�iB�uĳ.��֑`kɮ�+p�6B��C��������#�����w]��]�OA'�l�kΚ<�K/P�C��x�(�]Τ�8����J*8S՝�.Eǎ�.��*@%�42v�B�h�1��8?���On�@�K���v*�$Q��7W��{t~��qt�\�ơ�~���<����3��������M�A[����%u��=��Ǽ��2E|L���'�D}�xZ��	׽gK�}[&�h]@I߾��:��aGtx��x�Z/m�_O�>L\�(V5�g���"�2�9>����I"(:��h�� h���Q�zr�$�z��Lg���VL�n�Ox�tgޙ�k��e��,��;"\�⠁�4Mhl�?���M���OrB��:�e���f�/;���>a�=xz4|�%:�P�N�F�����+���'mu^�]jZlYO�*��/o���H7T��iAY�d�rޥ/k�VZT�|�N&�$9y���Ԟ����m���y�	���AJ�Z%�\�(~x\]X�����l��T�6:�k�q��>:KIxߊ�[/{g���[��֮��}��(����m��	�`���|�]�eĬ�с��-E}�C	���`οy�sϑIP���}b
CE7j����<b������Wx"�\~�:�v̺ʐ �Y����Ż��"��ux��� �u�.�uN}��� �8�Q@]�,�㑾y,832����z��W�)��gb�g�A[;�ʚ2���O�z���ʸP)��ZƓ�~	Y]O�B<6�P���>�\˘�xkI^X���Y�`�;�K�Y	�P
����04L-Z�O_k.ܵb��w`H;˕�5
,2��R[?�~�̾��cۇ^WyC�:[�8sy_,IVD�C�Ҋ`2�F��{\P�̪n��T�Q�"��sӺ����zT�G.�w��`}��_���֫�@o��d�	�6;��و��0+�0�Csx��`
�*5P��ł�,�;��y�v֋;��IRUOM�|��1���|�����JyHG�N{�k�Y0�td��q=وÖ�)�Y��:}���{����k���XOD�W��o#������X��Bu�y��6f^��𣲋ǚǋ�U@l-V�w+2Hn͑�տ���zt{�2���F�# �Q��;ZP�X�(��]Τd�\p�B�,��8,C�y"�;{&��?��@��$�g��њq�/��L3����C��Yu�O��.���w�L�3�ӬҐa�!ǅg��І���ڃ��l'�zm�RH`�i:"� p��_*��n"��o�R[E��h�P�;b�<d��ϠR��3þ��5�ӊ ��ue�g����������	Li��D��#��Q����6��;(��Nf�D�r���!�)R M�S�8��h_��ޫ�������8��-���^ܥ�F�;�}�t��|K���ſv�$�3�d��XG1�a�I{Zd)K1����y�A�/g$���>����s�и6-��1�G�)���Q�R���0-�3���d�.�Pvz�?���f�3�d��s����li��t�mJ�M��D�w��YS��{�W���0��b�Ӆ�,�p��M�$�>Ă�U����8�e�x��!��r�����wHm�'�g45&/d&2A-�;
���[z���BԥUiM<��Ҹ��m�:F�f,�=��x�W��%BY]�;���rc�ﲪ�k^�a�c�����õ_V����Ϣ�}�/��o�J�j�Qܾ�4(�W �`��Z�)�x��;ퟵ�C��@�3�����rG%�P˱/bﶬ�χ�Fw���)�]��,D*Qp��f�8ꔔ>�3�3�D�^Í�HP�Ckߒw�߮������������l�/��u�Œ�չq�����c�% RD��EV�Ja�U�j�A+K#L!�#g�*�y7��Ԉ���8�ȅ�el�	z���}�Sl�x�. �"X6FnC�N n��N>3۵C��2�)uCq6���^^�2��N|�.�2]��$����qn�?9<���g��J�1��0=�a2��2	4]��}c�ĐhH���0�1���#��rE,�����_2n� Y�V��޾
]Ģm@����[����fF0؊ڴfpp�[������V�=�Ƥ����"~F��ħ���Ik����;�ci앖+�l3�##Q(��F�eO��x�,��p�6 ��@H�+�~V��� z�֦����<S5(������6��G`vZ��DUYȀ0�{�`Gp�(#F��.�}��Y�2����A�.�Q'*���Qkq��O���w�Ykl���y�K��� ���%F���8�	s��L�@7
�����쮄�LL�$��^S��@�V,��J��#�����RJ�^�0g�#���:�,���'	�S65>���V�7��t��w�H�@f5;1�dx!�*�|�a�N��S;���\I#��%��k�Q��@yU���NJ@ۗď�nA�,j�����f<r?�W�|\����zܩl~ 0��0I�4���k�S�>͍�4݆ �`�,4�����8�(��2}��ِr����xn;�]8����N[�I�AA��cH��?U\�����T��lPwa����Z����h
����C�7!�o�	#N^�<1O�^郧u㝇KC���#25uפ���pż$�-��aV���;+4S$_���E��Y��G�|q�o��鈖��ķ�<�9�;��D:�]�Ũ��T��C�90-��*�)՜t��g߬��Nf�s���#qDAq�q�n��y�Q�Z	�u��_��C�A=W�_��wY�9�I��HYzp�z`es���t��!�m6A��-ޔ����h�T���d�P��_g�=�~��Ȓ�J֥�Kv���*�C��1�-�������BʜQ�C_D0>�R����%�����-DRû�B�t��3 .�r2��v�`z��� ܇�+�]C��YBiV�D�q��7�?�@-�Yq�e{5N84�]���ߞ%5Rz�$}�^�Z	�s��*��P�RN�+P�V�~� .�.Ś��ƈTi9Wg<�n-���"��� ���-@E�Q���K0�~�K�o��UƼ���ѫ����3��(��[d��"� �J�D��y=fP;�|�/��NHu5LkjwItMV�����VM�Tb�\�V3�;vD?0�k ��s,wR�L����e{\�}���w��"�F���j~�Ca�t��~ſy��*���	ܾ��?�J={��llX�Q�Ū��ޏj;E)Pi� �ua"� g2��~޹\��hEQ�I�� [���/�t#c@�y#c�9 /�cy��h$�5�����}5��V~9����'���K���-�fK ˢ�� o���W�F�N�{ۡ�,��z��A�I�y��gt�������4y����)�����eڹX.&��xb��R��o'5��GO����
a�a�D���"�P-��
i� �g�(1�0w���)��%�/�w�
��S7	Q��_�/8o�v���7R�!���֯(D=��%)�� s��,�L��Z��ʙ�l�r_�k�Ց6�KI^�JZY��J�X��_�G9#k0����@Li����tDw|c�m�*���K�̒"(��.�2�Y�z�~�����@�ש�R��2�C���;]��w���kC{����v���"��S�$�ɹ�������7r+�	�0c^��4G=�o���Y����i��F�pv3������L�Ion8i؀��&#BP��\T+DC_<�+�J��3#��7t)���>F��m�����$�YÏ�M�f��E���0�]��O�5H���	~�օ4F$��� NN4;p� �[�x++PZ���=��}}�p�a˞�X�,$�CϤ�����
����75эce�M�]SN��ϲ��;�.��YC�R������tT�V2s_(���9sh"�c�yl�U7JviN�FM-{����c �O�8��1��^�mj��a��e�����J�h%�[�o��B3��:*�~�Ծ�����FhỪ<��u�l�)@j�Kk����Mm�Y��]H$�Bf_�y��6�5�Ц�t�xOO:ȸx�/�"w O�R-�A~Jv�^2�j*fo�1�g.p�p����VKǫK�#�X��$�{_������3!�����ʖ6]�ʼ<�����$f�@��u{���pn��"�^O�h��O�}�������ڥ����6n�����~J�a^/�����Y�i��g��������Bv��S�M(ҧ�00`����h�r'������2���h����nHl�s�.k�z,�}��6��Fl�D�v�!��3v�նJC�w� �ߐ��-��fb�l�ݻ˟Vʝ>O8i�%����&���*���_�~��_6Ow�_�!tO��$"����Ð��&�����pi8���m�0Ŭ&ji63��to�%/�� n��o����t3"_#d0A!Rfw�x��:,
N������#�E;�5������_�u- QT���χV���LXT�ڦ_׸t� 2����c&���������f�; �w[��j�O�����N*Ǚ�Q.�A�o��Qrn�y�0�jA�'pg���/'�\0[ғR�g�&�8-R���Q�BR�L���9�0�j*�R��j�		��4#"?|�"QR<Hĥ�N;�!�u��,������9�n��C�I޸ܯ�E�%b�e�/��;㚑�'���@8�,���y�ܑ=��0�Kޙ�Kw��#AE�o�
=�^��\��N��#�<��K��������ЍB8d�k�ī#���.�bCE��?�>ccfu�^V�_ulD��T�+2�'�!��� ���[�b��dξ%�n�VNߠ�\���|^�0�M�ܔ�6�m,���U��F7��8�sn�0��K��I�\��?y��K9��Nx�8$���:��³��_���#��_3��P�E"8g�~�m2C����WC� #52dɓKq>�Y5YԔ(�"�Iu���H��u̵�ߜq<:�g��&��6���ۯg�}~�lDcT�n��Q-�iV��_|"�+Vy�������4�"]?~t�w�1+
�� ����^��	�Ln��<��i��>͂��"/J+;$�M����8���Ŀ�Ɠ�\���\��`aXr��tO�]�%*׽�敥ʿ��WhY�Ũ�\�	¨ ��P�IU�Ŷ�bH� ����=�Xv�7�ć��Hx�d}�/��3�����O��*B�G�7�w�NIŚ^<�$��1>�S��%_�6 E
�x��6;��/`¡@���#J����D��?���&ʵE�s�9dXT��B᪥2*`�-�S��7��Z�H?'�(����6/#)�w֥U92MQ�(���Xa��-��
[MY�G���N�kR��9��-!��K#��B�{{M{v��cq2b�b��>�ºmh��ڦ�?.�ׅw��d�dp��g]�Bu4<�MP��?�m8i9>&�����q/ϡՋ12e���Kb��x�p�g�nlt�%�ƀ���{Ik�:=�ӉY�����8���M�YDb�w'H�E�@��9j%�g�[�c��!�@�_���vʟ[����7\<�Dr	n���Y!���i�
OD,���U���֧<xɬ�o7Mw��L����Es���i��$A��W��7����V��s���D��Y��2�L�W5ݨغ� eS�NB҉���6ה��̬�.���u#
�N�0��y)=H��,1��g����wDe�;�~|^��u�_L�ґY�h K7)�g"VM�l��Z6�V�/�.�ɑ��Ϭ�$�n�P�{�Y�۲J�*Sy1	�-���b'����g�p)s[L1ۧ�m���m5Fpܸe��!6�D�Ѐ|�c1���Y8��'"���VE�q�8����U쾩�.�,BKm����:�]��ޞ�Ցh�`�����p�r���8/���y���i7	I��b�#�Ҝ.��5ouAo8+�VPWG��L��� /�P�U2XRI�jW=�����[j(��,��5�2�p٦#�OI9�*��nS �ٙ%X �W2ޱ�3��_��W�ug+o@��x�� ��a�8I'�*7�\�d�llr�Ub�ަ�@��0�B
V�Ӻ�.���v�t����X����`�M�m����  $ �T6� J��ȣ ���!o���hP:bL�Zf	S��A~�n.�X���#��l��=u�����H�	zN���%�����M,�D�:�yݔ��VNb�%�T�JNۻ���da�ӈ;�\<551,�g�au��g�jk��&n��Bd,�L��"k��:��MsJ�f�bB�Ju�U �"�3¾�)�5��	���'���V��(����o����Ȟ��9`�܆+T���j4�8[.��R���㧑)w��c]C5��G�����C�r)�v��9D �����m">R�kQ�,4{�84R9���衡6x)�-tJ�	U�M��^�^������u!���-9���u�0�1)�� >�>�-x6d(���l�ISp`���e_��\B��G��Pn����+7d�l($�+;������?z>���#��������	�?�¤�G=�(�9�fQ7�Q��_2�C�
"�C�)T���S�x����h���?��E|�u�z|�21�����.3I�u���F0���sB�z�����O2#�����3w[�ա!���P(��26��`i�zb�s�go��E� ���tw��ĦN�]�h�V����Y4Oz�`9�(��y�PyZ(ޒQ؃81���=�x�s�������E+�D�����h�.�F.oq���������>�w��:u�T���F�I�^�#m���8��K��R��nL ��}��q����±|�o�*�t���f��31������\�9���ϋQh؉qR�
��?��B�Dp�T��2�¶�^�B����0 �j�n����;�����Uƿ����}w���!����}��&Dx��og�Y�q���ݔズ��V¯��j�i��SQ��}!`�3y]���G73v�B*��� 6�T��}�� ��8��I\���]�:6��tb�0r�qH�~�X'����̾,���cd$p�'�-L��I�1r�5�ޱ;�TS� ���*��ͮe��6�4��"��
n�w��	��l'|��y��7s��Nl��d�Κ�C�:�;���@�eT���!�>Ӷ	�H�y(�S3��`?H#o�)����X�wg��O]}+�l�$24��I�Dt+��E�LI�ˇ��C�Q��!��˦������Ce���HB�i�׹�9<�b`�^����
���n�k����,bNי�%i-��5���:�����ϽO���o�x_�i��;�Z�B�h>�<!����h�E
�O��q����c�gf�����L?���)��I�������c�C%:E</���1�Yэ[7P�U���7�ݸǵT����d���l,����6�&ۗ��GJ�7�������y�=�.PV�Qz.��eL����'�<�5��aj?As4~�Y�[�;�GV����<�m����S��	~�̍)�5�=�8��?�B��l�ע��D����4*�t����-��%�����`+3vI��8$�Y�Lbz#�v��&�C&�oD�E�`S�A���*��'x��v;��lw^�������K�cC���ib�$����j��↛�0r��~h�Z�(��P��9?�W��U~J�g磬鄯U4��S�?*���3�̶����	���=�z�Gg��!�7/��*�>��z�0M*;��Vr#S-�x6���l��~nݞH���u���p���yU�/;��Qׯ� �E�2�CE ��B(��p��%:��BE��5��X�?�nX;���S^؀��q��O�˱S�vL���x����)~��At"��F˅���	:� e�?E�R4J�����yVO�ƥs�o싛M��}!HhT�/��8�Lᇍ�-�w%��j�+ ��~]972��K��ܚ��uf����BD+��M��0ߘv�����l�9�977���p�����rx=A�m�!�0jcņ#E� ��z�J潴�2�F��İ�!�ذ���)j��If��=��m!,/ehb/6�16��{_��5�:,>I�ӕ~�c�y��)hʢ��5��Qh}K߲sD�SB ��È��ns^�\A�c��+�" �����+ ���k��Jҭ��v1c��t9$[,�b}=/�Zx�W� V����G����D���}���t<��F�[mbro��f�g�����JTK�;�d��Ød�[�Q|�72����$���k�HN��Nq�ֻ�Ȓ�n��˺�����;�3R��I]*�����N�����Bs�=�Ws@���n����V�}�	o��b���ҵT���u�-�)Ȣ�1c��jq?����GtdQ���l�&ɭG�H���r^����XO�/{֗�\� �uW[��� f�lcFv��:] �0��n���lM=~�� ���S{�"1�Ey1]����Y�]��6��#�u�;��	Д�m��
F�r~˱\�|'�m���o���!�����{�HV�g����ʗ"�?%�2���[�[�:����(;E��#hx�9`{��N���L�4!mNL��ʚ��ѷ���p���}�cn�C�@_��]����K�v�e:�q����S�Uy~�O��/�,�u&�W�*�.�f�|�H�.!1ڷ��j볹	�s�����ਔ��A!�Q�#WX�Q�I�>0��
�Ń��[��h��B��G�i$8)q�v�<�� �[���W���;f;y�=|d��H�Ⱦ������ߥ�r���{";��1����ɍZ$�;/��k�M��4
�5����\�Fr�|�iN��Q�1�Di��yo`�7N��Iִ(�}��r�"�Pхj�T����k�1>���)�5
�@�Xc�ǫ2B�_�tJ}C_�.��Ҥ#���i�N�l�-I\o� ��b?2�y��a@%��3[ @"V�Is˅���Y�#��3(M���Ί��o��#ǋ�x��?�|�;�sM�����;�\�� n��Cԁ�0,����b
��Ҏ�K]p��)3�2��|�~��fw:�{p� .Y�Db$J�����MYb�I=����/�`��R�Q��Lv�rev
��-����1"D㯺�.�|2�) �<T��	���N�2 �Q֒HV��9�����UmccP�0i��S�ߐZn� �cOC� C�Z��;{����eU��}@��can
\����Xx��yW�2�m�߿Xa4��6$r�{����w�Aڦ���)r��0ؾo�Թ:��
�ry"�nL(NU1bX��%G�����f(�0 �YT�@�,�����Vk��C�ѝ�tI|v��X�6��_��s�1\3� ��6di�hPwc=r�����~Yr���=}��T��jϗ� �\���a43��|t��s�a��WNHŇA?`mC"�0K��J��H\Mbl�P��?���8�<s/;i	��:7�~@T�3~����V���h��Ο�^$ke{&�29�)sNq2����S_�v�j�RK�#�Yzg7ZO:ɦ,���Dd��H"���Yw9�ӻ�{���|�P�| ��)��Z�E̓��xa�FF@N5{�����^)��G�y�ěV>O���f�,|�Σ%���|s�����NB���@�}��>��q}�њ*J�%����AS�BB�
��WZ?o��v+���Igߖ�����z����w��"�������޷W?��}Q)[?z������]���6{���]7�?Z���ea��r��k<������ϕ����yh�u��4�2Juؤǿ\b�BY	K�#��=��;0������U�AS�D��1�(�S�DͫRŴ$$;���3P0/�ݢ�S�+��*�J8�Ԝ�x:4�fCvq��l�k���g�D���@��piLYu{�lR4��g2h�z�O���������|�3�E5�x?��0��)���O��wT�����b�)p+Y������]H�^ݩ� G������+�� D\���ӮE'�Q%�S)���|>�M�.5b(�K���M`>L�Bc�b�+f�ѡ�OڙB/+wr���� ���^mu�j�p��O�"7x:c�����`�ao_r�r�3�Uvh�[.2� �<7�~��o��t���q��A���o"t�i�;�3�!�EiE�,4�qp? �\w��Z=5�ޘ��pJF72�{=&��N׽�H�c���MG�q�詻��i�����>�s���������΃� �P�%-�iM�|��zaa�<�-� A7)�YҠ_���3Z/f�R����5�U�'�
/OS��G���Ow﷌�p�������b�����
������v? ,O�$}}��[
,��q7?L��*��K�)w��eA���6�',@����? � ��M:aZH�?���Q�ڌ�֊�2�b���2ǒ� nm�8�������*�.�р6z��מ�-�����{xe�A�[f_�П-JX�9����h�h����F���9� �Ԇ� c̶Ojj+v?����l�̝�緼�gt��h=rf����n�I�V��D�i��4��de\���[I�[�yY .x�-��@��_Ą0��R9J�@֢Ý�B�Ӟ_�ʕ�a|����-I4���;�8�M*d`��5k1E�\fZҍሥ�ЕT��ftz\r�A�/��Y�b�����8�I	���fi/�й�e+Y_�c�&uáf�b��>�Gr�*����5�Y2�g�����4�ş0��/U�p �F����#$ً��2n�V�g���?.�d]hWlm]")�?r}ZL��hx�����K�)I �Ӎ�"˪� f���@����n��f� ��]n�|�e@
Ev�Ǣ>u��\cܩ�-d�Ӂ��$2#RUH�j���c3����~ft��"4H��F�T��W��NX�*���
W�>���Mz�&�߽��}8VW���{���)rTyhXw4a��W�\��Y䩙ڴ���l6�b.vE["�q�kGN�޾d�v�w�7�G��+��B?e"�^UDd�f��n>����lV����V��ϟ�x��L�Ȝ�v(R�v���БI��u$��D�{\��<��n�f��>��}06�k(�{ص��f�+�YO	q���,�F�B��T�%��ogc�R��Y�0�g�or�H�!Z��g��\̙՛�O��:�m�h��<ܒu��q���5��C�$�ŭ����qS����:����C}%���,��3� �6��2�՟g��P+i���X�|Xz�c�$=�t=��Qt(Rx�|�_a�\�5,�뢉�O���D?�-�b�WR%D�gk��su���ۉ�ls��.wD��:o�1�H���K��\�5�\��k�`�1�,�>^"��E�� ��ۥ���-�[�-> ,@ٞ�m��~�Y�ʚ��O��xF��g�f�6�[�*�)��0S��'p=��Ӆ��13b30�/������R"ъ�t�:���>�Vّ0�;�E�v�4��L�JC����R���"�q3 ������H5d�ɞ[-��l�&��Z��Ȼ-��z~��2��/�5�l��"�\b������+�"�rnͤ}NO���2�[s�^Rº�g�����)�Q90�ִ��#f
vs�2[��C�鏔fIJ̸f���,�f:��@�%H�bC��M$�$צr�=�y�˯U�r<��EW(;�/��"�{z�����{��ls���ށ䴊�g/Lg$�`��ͬ�(�̂���%(Љ��ٳ=�xz�|#�m�R��7ŗю^=K^^LKe��-����yS+�85W�d�^�J�Cz-�N��/)s��RQ;�퍍ـ�o����?����}�a�n.�����K�H�!�)h�/����f�=�R1U�	4;�t �|#e�X�)��I�M��rW��e~𹵬����a��(���#w����'/���ݬ$��<���Ɏ%N�L��^����i.ћ=f���c*C�8Y���un�ۿ����A��d�A�X�A���)p���;�Zh0�ι�d��`��L��c���N����:f�V<���<�Nנ�/��O��.��:�}$���<_�)1�Հ��n��e�j�3��-p���w{��Db���,k��̊j!�\�nk��2%1�-x�_�=��� ^冧��~��(�G|��[k_*�Ah�|��=�����Ѭ�*�!UлN ����$�(���]��mbTj2Qn�t��h ����&�&����Y�`�C߾,�sl�ٴ�}ba��h0�Y���ˑ5��X-�4���ojb�Do��c���ʸ���>At݅F��`_eه���sS��Z��^��h<ͱ����WR����3����f�Ȱr2Rm-C�:#M�UO�r�yBhP\�#c�-�VU�64b�V�X��ׄI0!�����`Q(��@�#H�J?~���X�`�(�`xƻ��a���D�Ar�́��ŧ���� 80��%����[����_�����̫ErH:�jl4�\L�鈩G8��g��۩l�hX��, �=	��������9��u�M���������=�
�]'n}�Ԯ1��5vND�������$_�Q��G{��B��zܕn�X>Y��0�}�z�4��"�Q,%�������U�t
e�͉Y(�=s"�䫑Ǻ�].�Q@�֢�{%jϐR�F�],��B�� -�#xhCТ��RQ��
��JK��
�3\���Q��"�@��^)���3�f�^pM�EF�4�P�U�`[�!�xT��$(�}�R�KcZ�҆�bQ���[�m��h��3O��flvy�zh�j�?)rnY��Q��m�nR�t��y�� �4c��>�����0��
�]3�����㈮h�Ԑ��P�!z4)5a��S�/sa��k[铣���@ ��Qa�2Re�5͓����%�=�st���C�hX�wG	����v�:��D�g�bj�n&�i�xm�ob�n�����n��H�@��Y#��ۅ��$� ��|S�K'x�k��-6�p��و^���}��<�:伆?��8��B��Cq��ib��q�����Q����{�=���؅���M�z7	,<�Z����֥/�.I&W��O�q����8zð��E�:.��.�S>9F�]�AF6�c_����UVc>���$���#
�]3���)��N��Y���{��1���L,;~�i1�^��e'W;�5;s����j�qaO�a��$��}�S{𻳢�y._��k�����vqGL�"��.�X�o&�>�uU0�,,I�Tၼ0��	��= ve�r����Ľ5D���}=z�/�_�����A��|%��3o�"�uXbλ�hܴ���i��q���}Ҥ��{����Aȡ�g�,�d��J��L��/�]��f�@ "�C��٧wB����?t|�z`K,c��Gۦ����lj�g��3�o��'Y���)�)�:%Jwy9Wh���o�q?|1�m�G�5�
�1-m(�D�7� j�y�lLOJ������ON��vL�@�w��b����|�2,�����*���ޠ��* �.l������������z? �y
wM�$�E�)��)@��v��ۘ�Lm��v�"�����L�;J+2Εˠ��,e@��e���
��M-��Lfɂ�%(�Y7F�|j�~��m7q�ťOBz/�[�Q19Ư0gd�ס��g�力���'�+��5c�U���W�ǰ�o���0ƨ��������LwSA�P�Z��ܟ�!U.�����͇V�Y��}R�9�3亮��,/ ��p�ϑ?(�����`a�/C��	�Y��g˗���F��m�[|zs��ʎ1��p[���A��G�:zK�-Ȣ��+d�{Ew��q-��ʫ�lb�R��ޯ�J�k��[t�:�qB-X�7`B��#]�1��c'�s�F��ŭ��~O�C�7�e��I�Spy;�dZ��l�hW.A3�K#\	�4��iJܸ�w�pβfg��(���E��s�Z��1^I�����{����k�ЍaI Q�K�i��v�ŧ1�хH;���tȉ��g�bW�f�i��e
�i}��+]6ckz���[b7������,�-��~<N�`�ntw��� ��`��ڔ4}ϭ�~��m��=�VS}����Qb��b:�^�SV�Jdc*�MF��d�W�$�J'Kj��9�v��H�^�w���pY�$1��E=�\*Y����q7=��|~�G;� �e�x��i'�j:Ý= �`Qz���b���^�x���x��҉_�B϶'���Y�����*nh������]7��Ĵ�\¦8�cpϬ�u62-�Po��@z����a%G*D�9���4�U�� l�mi���f/�j$�3>}I��ڮ.+�!�Mt2����F� ��O��ağIL�d��T�q�&�Q�/��	F��j���I�vLR���
�F��5�S#�`2闢Q������?���O&�][^רm��f�9s��Rh�ɺ��>��\��uL��b�W���[Z�]y\��5��x졲����BO�������B�RMOd��E�3׫���KWo�ww�j�l��د��Ꚙ��
��(ǫ���6���;y�@҆��[MIPİn��S����A���F�=��Bd���v�qAc�6}�a׃e�3W��~�c�!�)�
�?\A�D�eo���\�4���tg�gD׌���D\a(���Z����������4����X��ˮL���KƋ�>��l�qs���Zd�1�Y8�S����ӹ�If	�ݼ+�O���3A��/9Bh�����������+�^�ٟp��^j��:�90I2���3���.~�����0%�T��}d�>��ӏ�,�$�i����8Ö�m��W��	4�CS��::7"Rew[D�[����[��{�@�!3 <��6f��bfF/%O�� E%�%^cL�u�
{�{�r�;���d��rE?���ViW}B�K�|��w+�G����>�1ګ�:���w���E�ڧ��?T��	Ol�h�^�&��mC���s�N�nض�O1���7/��d��D�TFS7��뒥�r���+S!���C\�����)��1&��i��:���x�9V�����	n+
�MI��?)u3����CWx�sN�n�5I����Y��[0�����;p�Z��s�ʅ ��:��JJ������6��zO��+�Oh���������FJథM���s�7;�Z�Ӗ��"x��f6
M,�#�Yc�7�C� �VM�-������$OuUs�^�ɹ�)�ziܙ�\��G �"�3���f1π�[�T�½�G9Nc
!�}�l(�X�!���b��t��ͩ����Ȭnѭ[��:ͫ�NP�q�)�>jx��pي���+�C�N
������^�-)*2�z����-0�V	?(��A�Cbm���f��z_�����{��������o���L�ꗕ$��j|�r�<6N��ܠ̦�3��u�K��5|��Q��x�Oߤ�iG�?%q'��z��,QNM����@�k�*�k*�[�?�J�h,�����N�Y>Cm����(����ĥ�c�sAk2?�c�=��Cˮ���h����=:
f����u�_a����i��*]���HW���MU�C�#�g���0��c������/wH/n������{��D��k��	*���v��*хF\ރM]�`��,��L��H���Ku�z����?�Y4)Zn�tET�!�RH��4����B4c$��5�(5�����sU�p1�$��&JzH�Q�j���տ1�a*�,Z�I�ka��>M):�ΟaQp�R��3Y7k���z����'��8����`��� ��/����3k"qg���0�2W2��"��CY��5\H��)jS�QC��L�T�܅�{�7�����.�Ng���^����kfBLvԷq �]���V�%I}��9����3ށ�I,U\��{�0O�f�^�25O��yt��9�1q�M�32�{O��`>�ܟ�c�X@���Q<�"�-L]S���*a�M�q1�R��osb�>��w\�>����e �hY��`}��$��
�Q���y�˜��V7Rm�)��;��1��7M���s���3)rw"���7SQ����AheH���="�}�Q�Z[i�G�H�G�5ߛ�7�#�u�Y�(\��b�XW���Q�i����g;� �n%�WQ\��p-�g�oe
�����>��{F�wo�}ϩsd�:ڷ�R�?��vqJ˾������L?�m!_�};;���L�pm�TȞ����^�0����N�c�&�Hz�Sa��X�p}�����������9��6�04�x���I�C'G�;[VX���pyT�2t��5x'Yʚ_��f�m?�.�q��au)q����RH<�"�C�bkv�;?R��t���?}��Xqp	���� ��1�M&�Q�r�J�Ҵ��D�PM°�A?���O��l�$��1���>�����Y�]`����^�����H��j�>Z�}"���*(O�x�&�`jL"����n��ԑϣ�o`�P���x3H)p���H��qv����eӖ6���T���5�Dg"�!lC�5{2 _-/��>caQP�j��, �6�q.~��U/��H��>ϩɱ��|ćh�K��zJ����n�ص�����!�F#p�����+�?�Rp�>�]��~/z����$�5�k�?4i��P�A���Ksleu*��o�����!���X�￱���w��l��E�3�%Ic1-� ��t�_`:�����I����^R.^��FQ�/Y���[���^�f�����5�àٵ��x�~�����X�r.�$����̤�ն&aQPޞ۫��S��;�x��������u0�~k���&ӱ|����xXd�8��e��Bs��I�s���7[�3�����th7s��چx�x{���;�B�?9I�y��
(�����s5�-�^����zp>q�#,w�n}V�ѝY��@ye�����Z�1�|�9��!u�2�4���7s<��k4��_}0�.n�/���B�qsʩ�Uq��)_��=����c_"�s�U�K"q��-��&J ��W6�ʿ�(^F�3�8�`7y�p-Q��>y
��`��K�3h ����2Ǣ��O��<Rr�b�Dzk����׸��ڲ_M���A.�E���*}����v�C͞'�jc�2���X�ko�@rزWN���{"=:/����ߊ��V��l"?�l��l��Ʈ>-��d}5>�!г;����[`��n`�����ARG���5ڃ]σ��XI,�(�o_,���S��h̰�wL�}'�����C������%6��Ty��������<�������d�-�g�����E�u�/���Ϭ�w�B#����B��h��+ ��
�(L��oH�B~)����ww�f��r���0���)���{��\#��d�����=�w�X��1���S3�'���T�K��������H�3ַ�H�W329�1Mׁ,eb���S%�n��A3^�A �W*r�;�g�ڟ��ϧ���L�_��:ۃ����rc�]0v<�9��2��G���h�2���W|bT�����k_D� ���b�E0<���]K���ԓ��^�����s���	z����^�j@�`c��c۪��E�E�:v__y-�\A��*�"����Bp��AHx՟���#8���a��<H%��"���r��'��\�K0ئ\A����\�6y��,�����}����%��[��3�:�Q��=y�k�Œ�/,Iy���j�n�_����IZ$�N��B�C�eu�kО/&��Di-����\� J)�O�e��UO4g�J�P*�n'g��'e|5Bť���G!jUnNa��b�S�������P�y�)�l�c�>�_��
���dKλ�y0�_�y�5�Z�_��өs��.�pj����ܣ��Y�+;+jz�{l���o�Ѿ��e!���6ΐ%t��Bz��iN^|({Q�v�z�[(h���!��P$0��Uf�rx�
����"�BT��|G����N�-G��˵�7D��_��C.6z�wq��� EP�i�io�0���ic;�:@8>J�b��&�*�9u����t�Hñԃ:/a�f�Z��Zr8ɴ:�M@�S�����УY��cy_E�\_h�8��	b��!C���$C��b���<͢�p�-+�4�C�%p��C�D��Ұ�����M+��o`��p��&~��eU2�cy�<w|���t�e�!�g��ksbʍ!� ���P��h�ڪp��1�6�Z�y��9�-?+h�K���x-S$tp��I}B<�\7�9*�R�dsK����WI�tv(��`���Q
��g�[_�m�~|�&�\ǃ���R[֕��x��j�gN��$��o�����~
%�k��a�s����`��X#�����t���t�����N?�v���4���͙٩�C��|�@�QyEPJ3����h�e���i�ov���+'��<�10Kl�SqM�r�v3b�Z�濸��A��6�ΤCڷDh�#96 �����p�+S:�{��|鹅Sj�4]�,���`���ER�rq���$����?k1����{lшn0����pn0 ̾}��8M�ɞq#~�oq�P�٘�Nj������w�ZY¸��nh��n��x�ͣs��-y�Pi��y ��lv�RY5:����p)[��W�SV�C��|vD������j����^���v-N�W��A��Ӟ]uƄп���;�K&ƺ�!zJ]����]���.��,w��da�*�H��O����weX��r��ERN|4g�h]�Eĥ|fUoxz���.34ų�7{{y�7l��D߆�\�X�5��zGj��W9��Mwp���PV�P�m�vJ����� nw�~1]�����.�
�P��S�2*�¯^"bI۔H%z��,�?$�ᴷH�bS�>��d�Q
��l�a1c1�H\����������{C�����T{�%�z��5��_dD�G�C�7�U�T#���{�)�K��̧T&�*�g���ڒ�Hw^�P�i����¥����z�+��S��,S���3��]У���h��dJd�
��V��eΠ⯬FGҾ�����A��Պab���7�r2���U�[�˳.�t�;�WC�h�ɀn�T=�[�1�Q҆�p�U������
Jv�}F'�{|?���2*c�JW���}�W��I¨�������b~B	lo9,_��TƓJ��7���ig:P�7�P�����j�%�\;l����K0�V�M9�Szϋ�~����`S��3����]
')�iK��L2�3���G-֨*�LkF��9'8��
�2��g���4�u�#3dpC�j�~�����b��:���	�jO~O� !:z�p�}VQ��̖�������D35�� e=I���b���}X�k�	�����_aA�����1�9�	ѴR�f�q�<��&�ϣ8etHm�)�7 �?M��dҩB�27M��|�9�!Օ�P��P���	�|Ѽ����ٕ�ᘛ�N�&���x	�w^x�4����U��{@M,�^͚�j���J��ݏ��������H;��[I������-�U�ݣ@�H��-�ڐ�����`�����G�q��GrR��A흷�9�I� ���v!�fz�)��'�&V���`?�}˾)�%~B|F5%4c��U]h��5ǜ�����@��1p�m���>vý(�Q�(w%%�\*�LLu}�+3�������F�Xޤ�nSL�'�(��´�	ٱ9�|��3���D��N��Ĺb[�㏞ɽ�Q��QL!˿��].���t༱����*�X�帵�y(^�k��� �Sq�V��G�l��ˀ����PV&L��V8-ڽ0^������c��� ��3��-!��Ժ�j˃#p���h�|���Y4=�����@�*8gbS|��q!���E��D��H��,%��4�[a��4 ` `�0y
�dI����vP��S.Y�/����Q��M�X�% �0q�k�UD�Nn� Z����.�����S|\�.;�GU�,�F7�X�����C�Ż�5�z�O���m����	�z��z�V�j6��@$�gD���\���\��"��_�� ��Ҳ(RR��ϣɄw�����[�R�,�� )�xO�R�P�

�Ghd-;|�2v]��ýV֝C���2�\|�IWF�#��k%!VP���|Fz�b<��u�pc0·jv��#ܕ�\��i�ZC�9z�
TͪL"�<� Ӌ
�z�����x��;�Xz�����M�m�I]���4��NiF�qHD׸e[�%Պ��$��_ڗ�0p��]�8��Bx�(jȹ�)?�� ���<����,	L�c3 �x�:��!܁/�݌��=����+�[V5����%l�� aI��K?��#a�ּQ�Z�*H?����)�EL���Ɓ����6��%f���K*p���U�����pc�`	:���:9����%�S]���488=����xCxvP��<tJ3�j{��|-�7N�8� ?���܈&P�bG�;z�s����n0�U�j���3���&.���� �k|_!tۿ�#EwHp^�V�U���5��T��Y�96P2�e~Z̊-@^ֿ�EK�yx�2�l����¡��C��9��ꐫ|z�����Ș�ْN�e�:&h	��۱�/q��g�}�ԆH�i=	�;�ғk��63�xg�;�#�PsOq�@�$=A%�O��$�<c���xa+hY>�<h��ⶦ�]��:�B3R28����׃��w:Au ��*�oa(��3�7�R�T�-^�߆�?� M�OPP�
����d���$jz�X�e���$G�?�O�Y�|����!%?�'b���ٞ{.e��`��.W���L"�fڹ�S���(��5k�����;�0�
�Y�q/������6�,�N0E������QP��H��������)�VȭA���Bg�³�P|k��T%��s��%��V�ۼlZÖofaq^�}R�]2u��]�1�h(��N��4�3`�e��QU,M%��&������R��GJP��"���wL1�&FV�H�,?\���v��H+�Q0��.���� �����+aV����N�۾u��h�����$�sALH�,�s������S��ocx#��j�W�է�(��X[j'�_�/.���z��yb<,�$�� *���U)c�z��du�>�K�7Q���W�JU��fZ�ٝA=j���|B#�1Fa�Ь��gy��b�D�^@�P���%cپ�j$��ΐt�`�Ja�������Jf�r!�o�,�*
���c��;�Ќ$��B�5�G�H�q�!��*m���Ր�H��T��w� H��P(��2�%�tC�|�,�N��\�>OI�>d��-�G�)��O������f���-�q+���2'��J�ܞ�1(��M.��f<$��T�X�|G�<u A�%D��B���B����R�*�'-\v�=e�`l��O@��W�򄜐���6�X��$�	� ��w����b6bܽΖuO��7��7�����h�`��-�`��E�Y��:u�=w������?�{�A쮱�,$�&e�T�A�����ǎ�2��F���k=&�2��7��Z�E��P\����,�/�e����!b�V�?��R#�����e���Ѐ��M}C
�������_�_����S.9�Q�*��1í�w�|���a�μ_�f�L7�T<���$��ۑ��r�9a���S���
���vr�T��vՌtVp���i������9�V:)��{,PQ�$B�,�jZU�\�xUqrkת���
�W��7Q����d��⪓u�<�+g����9e��И��y���������R�-��y��;�Z8nk����(eS#Z 0��>�L���>���ߴۘ��~���\��"�Ng����>���ػ�E$��9�_K��9��� �����9˫J���D�P�[�QE�w�!}t��.b��󛒩:c��`��5�O���㚕�N����6޾�?Z_�"8K�o4�0��Ӯہb��]��L��&��oX�=2�,�����'�4'�!�n��Hcz�څ�6������#o�-���׫\���z��^�+�M���.F;U��?^?Lr����ʶB�	�J����o���szu�CԎ�7�IIu��g��&!�6V2�z��ۡh<�����2�����|�Ϻ�c��w[���;�OP�mt�S�8c�4� _���<^�N��/���K�� hJY����%/�m��
�N���f���`�K�����cX����#�W<�*ȈG��vA4rbK*��A�`�_�	�����	�p����]K4��+�Ur�����,Z�����,w�� +hSY�Է	2���"��Ye�U�C�Z�Q]���7C����i��I�=����?�Dz�=;��7�he���]o���
�1ԉ��n@�(��!�X4�iU-����x�t$̝m����=��iv'k zL��4�������BR�;��D�cW�"ܐ��seO��T�uR�������Z�<��H����F��#p�h��f��0��[�L��Zn>�f��m>.J_��\bs&���hZ�jf�(Ga����tQ�����Ը�h���m���<�����y�����:MґW����c!5�jpN�肍��n��}��i�:tUx����+�7{䗇A��F����W��#iW�_�zkl�4�qz���=|�Ջ�T�!��y����
"��vgz rpT���������P���s��)Y��=�z�RU�#x�����g򙊯�"����\��Ȱԛ��sI�]����%Q��ڐq�;Z3��,����~�G��Ɗ���e��׬��yڞ����]�s�5�-4�%���
���}��6J	/V86��� �Q�ng薠4�.A'�.6��I�ù��Иc���gH��nZK
�lu�7�,��[��U�W$�L6�Ǚ&>��_�2�7:<�	c>Q�;�4m4/u"}�Z��O��S�6�M�B������,IQ�Tp�kL\P��P��)���:�H�{��v��{BGG �KF�[MQ%ڟ-waS`�i�-Fm���/JsB� %y���S�N&A\S�n�,r̲V(����O��&��YDP%!u�P�&��gJ^����әpt����<xS��HC{N��&�Y��W��P,%Ǟ��:ؐs_ ��KƎ��
^I��RUmT�~�uj�S�,s��9N��H��0_�%���60�}T�i��¢���{����o�Liv������Ɩ�EZ�\8\פּ�@�N�*�v@�Ȧ_���U7�ƉL�sÅ_�0�I[��"�𩴍��2K>`��Ԥ�H��ɥ��w��^�ب�ux���T>�b�`�q�Ⱦ�w����T>_�N�d�=(�\DҕL,�һ!��M <��OP����v�������{���ph�,�!W�h��Vhp��A ��{(_z ��$���+7���	��|��<G�?4���ڂ�*^@���P�����-/�\�"E�lƚ� �^��W��|�ⴰc}��W��4ʡ����/N�G#�����*��v�W$G���漥s�-K	+SX��ʪ3+ޅ����9ʲ(�M�3��1ڄ�El�+��q�k�zwg	��;�2��[}W{��s��K!@4��{M�7��o�s?�kc��؋���,9�2�"�.��>3-�p 6#��A[4��1N鳷�+����)�U��7yZ�?G[���m�\:��&\져U��Ғ�r-R]z�d6n��t��q;��:�Љjyfx�(�� �E��N.$���@ ���Y'��có
�fPQ`1:�@�ِS� ���a	@�q� @�:�QJ@4�y��
�J�GE5W��o�E�\@������]�M�E(�R�����F?��Mߵ�|r2�� ��y�����keGg�矮M��������֩��&���A�ޑ�IC��g-����U;1Rw�p��[�]��{��C�"|�f�u�T"C�7-fn]u]�-����-S5Ӕ�O��W:�"+��#V�lY8=�S�p�S$	D�'`��-�E��s�1]c�Lh���,?6�~N0����فT���z�:c����a�Ј�%!f�mG�{�
��9���.�2�n� z��<�4s�M��^v��+VҏH��h|�������s�=R��T��f�`L��$l��y���G�ژK�z�_5�R�n��h�V@�C)H�̖�5��G�@��D������#.e$T��+1FPb
f1��,�1���$1@�e=Ћ+U�r�+�h�3�ߏ ��t��8� z�\�>�ɰK��rs����,���"&�}��"���"p�вy�� H�p����
Wc���^��&�oɅ����ෝhg��.lk=I�Y�y���l��Q���b��W����z��0���R�� ��jn�J�&�
�ʽQ���s'�	zH�{0ӥ����2ѯr�n����z�ѷU�w�餧��<z�CU:�yy�4�(��4E�&�W��[�/�j+�jƋ���F6�������{a{��aR�XG�BG{y�(B��T8~��,�#���<`:� �m��r,Y+�$��'�׭Ԛ�Ԩ�����kO
gܤ�_+QIl��f%�Lm�u}U��0�ާm�C.���V傧�䷫@�ʨ���r�>0fs����d:K3P�����)i8X
o	7D>3[@@�}�%"4)ȵ�L���_�=&a�<�\A���}8͋��+8���پ|�m������-�z�r{�ݳ(�;�LA�Sk�3	u^vpo�>��Gm���(-5��t*��2��bU8�a;�\O�X\s���$���F��h&��;�O��a<�^m#~ö��e�$%`��Ry�[�8�HFA�u+����;K
Ҿ�����;o�O��8x�3�Ze��$�|�5�9���Oiy��A��N�ؤ�1A��_!������U�{7O����*�r|�@�{~�6���Ahp{�8�Ũ�:�qv7�7k$19p\��U;��۝�1���{g���,L��>_
�f�
Rb���L<�aa�@jU�����VnF	C3댿�	*�΋Y�תQy|0ڳ��YM��i.]�Uc��5�9�n���U�����m3�#^����G�{�ɍ�E?TqNI/���6�kM��Y�C���V�=��	����+��x�>MCd9a>	�a������F��k���Ex�SR@­��	2�#rZ֬�U�����.i�C���;j���_�܄�]X�R2҇�(I�;=�7�^5d�(�H�~�����^�?��B��R)��Hߟ~8Ǻ]?��꽥vJ���P����S�\��)Z&�	]Å�0��rxȂ=jen���9�n�3���~U��蝦1��Os��|��5�g}&�-�}Q��X�a��(�r��rT�$�'�C^�Q�*"�\j1�׃X�2��E��"��)�dw0�m�6o<��t����C�O�&��:�Q��>��N��:���2���i���E%̲�K�
DE.ڔeW������O�'>h([����g&�e1�����������Xy������΄i=�Ւ��a��z��xa��R]$�� W;vO�seE������j����ݍ�'�",=�=�m*��u��j�TktV�D醙�b�m��m	��AF�w_]���W`�D�B�g~�]�ˍ
��T= �8M9�@�Z��b�I��-E�O����K��R�o������;%����q����2lQ�-D>�0Ma.�y����u�)���#yP_��3��il�A�P<M��j�d��u�t�;�㛻������%k$��x�:#���u��/����i�5P�Qr�Iý��*��,64�;�c7g�jU�Kw(�if�/�3�&�������
	��x�h	�f썐r:|n�~�x�U��En�z܈�4�G&:ۏ��S�07�ET��!M���.'M�z��"�~Z�5OW �'#��m����A��v{>b��h����^L��*�O'�r��$1��_��
gl�#����8r{�9�-�6��Z�c&�&w�8�`Z��(Oӆ����3�ͩ�;=fG�g)��Ԓ�7w����0kp�)�N���J�KC������EKjN,B/�3�F���Jv-vl=�L�ܲ		H)���.���3�h�+�߁@�幪���6j�}�I���r��t�){8G�O�#U_�1��|Jb�4�8
���%�K�l~-C���� {YBݏ�{A��G�C!uK�䞧�&w�
-n�!�}i����]^��z����E�κ��|�V]�t� ��2��E������l��+�a�K�g���zĕ� ~��⪂���0b�Ww�C�Y2�i-G��H��6?�{�N����ݙ�DP��ƒK4Vh7>=m��j��6( �2�@��U��''�;Rv{Wf��[��W-@;�e�{��p��$��qxm
1��f�8��Ą���C��zZozeh�T@���q�ƻ�Ʊ�ͧ�LuI*H��|w#q�k]����δ��ha4}��ƞ+�v4���"k8�Rl7CS���H��4���\�i�����c��^V�7x��iZSh�f�+�|����a�D�z&��:�|0q��0��_�l;�]b�ӱ���}�z�W��G���^�!�h�S04b��6����W��Z��I*��=��H��}L�'N�AD`�$�Ё��X��_�{��y�%�Gq����!�_6�Omn��DUS�J܂Ζ��N��ԃ��ׂH��UȜ��FBd�;6oSe]�/1CJ֮uB���q�,��U���.�� �+O�;�%l1�X��}%*��˝��Xxt�N�5h�(��J���8k�D[�흹n�L�{���jgA�r��9����|ob��Au���#A9+��!�`�Ѽ��4��P���>!�@�9IP� ���w
�B�<#�`�J�RN�)��U?ŖhV�F��zO�ҹ�{`����PޕS��7&��Z��@{�:!�<4  �R߯���h	�����R���Z8:��d���?.�!"4��frxp�Թ�E�����
<�R��C�rHuM�rU+Sa���IѐzJ�r�oҬy�@�}A�����Ʋ���'���*w��ۍ�R�=@�Y\;���|>������l�ä�F�Ձ����j�Mg5���N��Q������  やL�6wD����pI^�e� ��M)i��Qw{0)8�+he�y��|�{ǀMX}��>�߯�ۉX��JW���
��2�5iɋ��87�h��t "�t*ԮH��&^Hg�7�*�p')>�c!s�����Y�T��<�J/�F�ɶDfڦ���SfS�ʦco9����x��G>N�S��&k6��p��7^����e��h�I�Q��g�E�=y����5F�j�W�(e��6���8�G�l<�j�j|��!`��o�S#,���lj�Q���_s��x��0Y�8���-�ϵ3!���T�=�,���n�6���`n旟6� \kZc�I-��� �p;��4��)�r���	��<�wA���F]s&Z�Q���M�����BN�c}��P���=AM`�!)�i�Jܜ��@g&��:�o#+�>yt�^&�.��n֪� ,Wq&��\��J�h��豇���j[�}��ARP���Ƞs��8�QiM�����	x�zB�?�"^C)U��U���!
�0$]�����5�@rf�EB�cT?Š�+]mr�ʣj1l�Z|�"�=�� �6y0Q���a��.	d4�3�b����)N�Y;{�<�Bm����J~�w�$γ ����c6DɌ�2%��/�5��r,��REs����7�:�aV��&':d�ϧ�u��N����[�/���f��Z���8�Q�c��B}gc�:�G����������B\��P(�F�?@�uJ���1�A��V'����K�#Ǔ�����&�`�t�n9Qfx�|�=���x�y5�"k��0��A2��a�8"`L��Bv��D�	�x'�eB�HaBhx<��A-y�/�bD��ʎ��ѓ���.�i~�����]S +���9�hِj�ƭ���ZۺW��^���M�#�s�	��ץ�Y�?��`ƶ��
lP�����-���j�3���P���0*i�c���ZR�I$������n6�M`=�Ϊ��Y���^3=i�C����/��U���`Ø�
!��@�6��(F�O<+�� C*�����1���/��54�~H�.R��Cᶄ?;�6H ��`��}�M>���:x�~1e@�V�:3��Ҁ��)�0�4T����o���H$��%r�>�2��*pqP�ft����z �.b���s��o6�Wݿ��!�$ 3�6L^�`�1��������|Q/�f)c�%6!�����kG�ʩ{@+�]R4�S\���Lߤ�5}�D�(�A#�EؿE-K��� �N�|v�v��I:�+��`n��u�V��qUN�V)^f��R�2~�gR&�|�8��#>�
V�L�w��!�<�Ѐ@E��_ü�T
��A�P\���T�fj��<�m��;��l��*�?N����JA]�S��/j,���e�͋�a�'�zS��~���ÑA�xMI�jJ9��@n5��Y��ʰ�ʪK���bm�3G�K�2ru���aS�鬝o�1�ɞ���pԴG�L煃S콰�JP˝���މ�*��?��3��Xo0$�pF��#��E����f��`&])�i|��?�$�o����9+(������i){,\���D\�����+��NE�6��69��*���qx�>��?2�4�@�8�0ReF�泌���ɭ4ᮍ��
�5�C�z�W��@�p�D�����nY�R�����Z9��U���}�ehP�{�n�m����yB���m��łqI'k6���ۖC@�dO��
3i@}�j��Y%l����˰����$�U+I6\���;��r՗�]I,�6���NͳA2�%�Zi� �)��0u�o���@u�LB?IO'	�"��aYLD��>�ش��*Q�a-{ùhjz�?`�����c��ܣ��K�m �H��a��">+|J��h*���]sbN�}�'��y@>b�C�n�Dq�<e,g�k@߽.-���C
�-�o���u5b��Z������
�#�i��a<��Psg��ӃO���f�����9��B��P����Ca[��#h�����$*��C�t�(��rP����XA������M�l,U�l��睸sg��j��Ht$!,BO�|��Z�ilS�h�x9���4� ��W$���Æj]ǯ?�u$]c���xC�f�gz���,r3O8c�7���Om���<v�*_t����J�=qW#P�+����A�k�km����G��\�xc^[�7����~�k��*�![�ٍ�p�I�W)0Y��.U�5�Z�7Skf7?n��j�1�Q^���6Ʋf��Ϛ��nQ�&L=�C�e�,:��jlބ#2��\C���}# �*1�a֔jf�o[�8�LtӪ)l3�tz*����T(bq2�A?����jrhq�ϲYLzcdN��7i.I�A�����c��g�z�y�螰���TH"�LҐ��H~��[1<���P�ZQ�ͫ���@ь�c�1�|y;¤j[�*!��\�q�]�6��N���(�A���0�=�9j��6�Q,�M�s��3O��5�n�G���X���j�(��7��#���ieLiJ:-㲂i�P8.,҉|�:��|��"0'���vf���ޝL�J(:��8Ê��%6tYRY�I��V�c���c��-F��U��~��2�=4���zW
5N;~��[��6��(�U�u���R[c�+$��qj��S�t�[<�~le�%4�ȡ��۵� ���� �xKK=��2@��jjCq��Cg8#C~0�a������j�C���L�7�J+w��w}r�G�i��8	�H� t�ad�y�3�!��>�J�_>}�}6��~��#<�Q�>�[K��Z�z��U�J��LT�f"����a���c�dD��������0����>��L��]*О�/�FO(��qM9���r��p�f:W,�U�d�LJ/�p��B��~�[�.qgt_�,$�&
2)])��d����ȹE���������X-�ƨ���O�=����7�\v�E��9r��'�|%@�d��]�Ҳ���SV{�m�R��rMҠ�A]�?�f�wv[�e�1%����e�sF:��,�'j{�Ä)�Sy���K���0�ʥ�&�ђd���Y�{�R��"׿k����᯺�"U�� /�d�Fƹ�odaɡ���r��������=�~	���;O�>ҴɅ��/���x�8�Ǵ��f�s�xr	R�^�)p����p��ݞ��c��qЫ_;��;�v����#a��"��9� 
z��Q�I�X_n���R��Ze�T�Kn��KO�c� �2���`y?ђ4	�W�����a6{<E9�ʎL��	<r/6ی�	v	<�n]�[8q�+2N`ѹ�<n�M,CJL!��C0�+7�r�?x�>v.!��Y���0�y�i��Y+��x喑��HL�:���A�9/[�}� 
8���?�:k��\�d,��2'������N�-VR��X�78x�<%%4��y��b�� l�4"��$�,�󰝹�Ȯ��^��`�4+�aX�����Yi�?L�x	�>�/wlQK������f��`��^i��l����T]�D��p��<ޠ�1��c���gIx_�;	m�5��B���"�����v��C�ɵQ��z�)5���*'�.��}���81�ˀ-3��	Cs��G�t/跋,h�^iy*Y� ��]��G����wx���2��@�.Y?�A�.��X'��5ݒftʩL�P��(|	�J��4)��4��؈�D(�h���|kEW�57�e�U��p݄\��x]�����o�ҿ��)y��v��#���z #�	/��K�,M5�����	����R�3�'|;�%7{���}U�HԧU��J��KQ�k�,�0zߦ���i���� �A2��t����L�F7������]gg% ?j�r�!�n��L�s�hM���K��D�ja{�������zUC�3J*W�4��Q�
ŒF��q��Z�t'�����h�x�SP�<Ib'�tg���5���B0W�q��?�]�_.��j���^}�[�&��ڀ�K�� t�/3 ��7�(��A'}Tb�����6\�$�B,;&Q'���a$hO��Ts_X@���/�/V�q#��(x3: I)/`?�]u_G~`�#��S�q9�lE��x�`l%��0���K�~N�^�6�-�U4t�W]`؛����[�2�0�V*��f���BO�8�b'U*ɵ�ܖѫ:n����*�
Q���ERmӗ_S�TXl	�^�29��#�^�r���l�Á|߰";�/���c���Gn�h>&͡��U(��A,��Cu�T*e�Y�d����J�nГ��F/{��3��I����k�?^��\m"�G���۶c����q��!F�V��R?��vV��p�|-w�"��8�r�o�� �|���Ȋ@�D�t�d����p5�����N���p5�^_�`,١H���mޟ�^S�ꄷ�ܴ/ٕ�B=�)�\���St˫ve�����R���݃�3��D�;W�@Y}yU�0&f���v��v��R����U틠L�	Ҹbp6�9�#��ȑ}}C�I1qG�WP<PAI���0��� V�`�"	���cI9w�)ݩ�s�#%��KC�J+�0�����v�<�%��3��4�J�!:�zmC�1gYg�/斑���l'�=JI���S�@y��t��'��0����d,����sT������N�l�*�"����hB��!�0I�E��������XW5�s�h���ˠ-��L�BV�Uθ�>?�"���[?���X�ߵ��S�pxKX�,2����y���d�|i��煜(f����W�H�V��Y ���W��T0R�K���E�?��^��Lw^���p̀6�1��{�v8�����S8V;��^W��������o�f��YcϒRR@A,od�\q�+���T��F�iB;�v�q�t��f��;<���B��}�yU��B+^�C���q/��C�8�`,T�Z��W;��Nwz�_� �����|�O6PT��(_�v�̷<��������\����A�΁��`d,�@���ί��!�A��"3hX[m\����o\]S!����Ptk�,�x�u��\�&=9�[��g4�@�$�?��?����w���l��r�%Eڻg�q6l�<�O��Y�Í!�Z�X�t����Pq?��lg$~�<�Q$n���*��/]��Y�h.�7���".8��*�=F0!��<t������/U��3˃�5��Q�usԨX��_<m�X������ꘛ��O�d��� �S�NF����S�9)�F��H��˫�OO���,�L3�ʾt�f4�����K��8��aS����i+E�S:��:H'Zu��s�B�,��������O]M���4�	��K*!�+�TC���e���U�$7�c�ZiJ��,d}�O�3r���C��S��J�|��ђ����_�����'8�v�
#�x���
5~##�8���LM�˞�tyǼ��eiAjT�t�qw0��,Xp(�{����6��R��a��6�-�V�Qg�ڨP�dv��84�-alQ���f ߫����x���/��(f�q�@�6���Q7�]b:�}�j ��W���9Su�e>=j'��[���J}�Q���:T�<~���з�7�0��%�a4*m}��ٯ:7uƗ� �ae���J��
FA��&W���ğL���-������蒅�?j�<�r-�����+�R��O�Wp�
�NҘ�Ö�)y�gj,x��M��}2���B���xu���9B� j�Rg��*��&�c�]H'7��,��2z�D�&�FU��7=.�9�z���'� J*{n�)�2̹!�"��"^骟�$r ;�t�.Z>w���Β�����d3�Os]� `�6��!����P���C�ɧ�\V�o����o����;/�k
��o��b�6�?�\S��q�#�ٛC�~���$�=y��E��[\�m(x���,�@���gj2�hY�Ήl����7ZƷ�S��_2�=ژW ހ܀V�}�[�JP��o��m�!��?g�o� ������Z��nr�Z��I"_�Wx�����l x�n³8ZN#i�s�L���T)�k5���Ol�+M��9�x�BT�_lCFu�Ķϱ8��֥w,�yxs��(�\(������MnA�uW���W��ךrv�ޗ/�j��8�hw|�fc�+�|�^�˽�'��Es<.�k�N�>O͗�/���W�'��3�uT|��'��	�m�Om� �q�h��x�$dE�-�;��� �����4˸����2d��7I?�U$i����O���a��5}%��%�Q��o�r8��>�� ���2p�����k]�Zm��6 ��|N?E;��r��{Y���Y�4>�ڼG���RiW����䫢�W��}Mގ��޾��}��+���I���	�X�U!.�D�#����De3����F���\���{���
AndT?�Ǻ�+�/��S�XX8r�m"�	��*P�Y9 ]�	-W�� r���Z�d���K�	R�u⑒᷃Ĝ�K�0\!1�����Uq���j��%ڊ��#5 �
.�G�ޮ!M��q&[�Q�(�W]���+�Vtɺ\ȑi���K�C�o{��S�e����ѐvX�o�#�xpB�ja�H��v��>>���cf�PN��lj����;��l�S�1k�!Ɲ�J(ׄސ�Oՠ3����3��IY+��O�nnAy��,[ޤ��z�ܨ`�Ț�9�ݩ�\� ��2�gi٤�>K	F�;'�^>
�]���F-_��f���g´%�/,s]p½XpH]�u�<���}�eC{S�D��#�M��C��@��Y`����nlt�����9�C��?y�Za)X�ei
�M�zF�Js��	�wu�E*��]�',r�bj�NB�1P�N�!Z
e����u#n;i#٫�u��<�H�*ysc�rRBt>� ��{x��Cj�pAŷ>i�����?����a�\��C�n����$�Z�ɱ$s��Zh��}����B���"u�y�x�m{v2��G��(0Z��(\:]������������ZXi�=�R=��B��M
��x*��tU��S�yŅ�� �����[�J	L/	�ކ��e��M��"B��j���|F/"�s=�
�P\iK�A��̨�nn@��O/��3~����mR��|aľ۹�d��W�8y��	s/MOR��~G'�nq{�	�
���ne���Xf����(�d{ٕ���H��~7�|���.o�u��!�1�Kڝ�+3��mͅ v�63�J��[㲳����A�u�M�9�v���:!���:z���C\ܚH��#��ݢB0��o�|v=g&��Ύ�m����ߧƉw��7� 7�I�e��čE��i��H���a��xF�QXB���m���
vS,��枟xJē���1SQ�'V����P
i������\���y�o��6	Oj �o	�[� ��x �h��>�0w}b󺀽u'���(W�m�,���L"� �ʑ�Oj8����_�x�g��F�v�-����tf�/�R<��r߉R����^����~���cc����ﬗ+lP�����ҭI�A��ƙ٩��̪%�����&7�����?N1?����ihZ
�%D������D�L�/:�I�?�r�.�d�ľ�[���xVe���qZ�E�af���,���c@�=�޸�9�1
1|ejc)��&f�h�Y��x8���=6B(�B�~Pre1�T5W/�reͅ�o�����������.Ȕ*����$f˿0}��܋bpE���ʬ�`���ǚO�(>"�!�F{���	S�
y�_Z�~-1fA��C؀���[)��E�-*�)5���U4��-'�,K�}TZ��9"��Kv~��)�����6=>�w�*�k}i����~�	�b)�z���ht����馠ՊkJ`�%�y��Rk�U�^���Ҥ��\W��wa���*x|Ĕ��v9���lL�,Esw����8Pm3��(!U^^ɑ4)bH�K �J��ё�e��/
��/��d�h�H���N&�t��<��v�ϸ�lR�'�d"w��
׃	?V�����̼���~�o3/���CSO����b�zWs��B2~�1�T����h�j�@� ;���׺��V�?LK��D�N;�"1��;�'�^]���e�C�G��`f�������Kg��� �H�[	�L8?w��
Hh�8���ml2W�AD~���i���ң�E��ax�K����_;�� ����K�%1���dd�/��TP���ȉ��Bj�06������dV�vo�����c��W�TO���]�*�B�3J��>;�HW����U�u��(J�B�+"S�ۉ^aR�4��w�a:�ѽ|�C�����P�z�/˿���QN��	2Zg*1SX����F6:<3+AH1K�����[p8���3cI7�x�OQa�����Ջ3�ږec�� ����oOK�1=7�F�����$d����1���~�rMk,�i��`�y�*�Տ�v�90k�!&w�O��|rڅ��K��GO�ֽ�D*��Ӳv��Ieȓ��f�}���T��B��C�!�un�H��!���P�՝&bЛzm�Tr'��}��o7냱el3��O��Wb݋u��}Գ^q'�}RD���a c(��������s��*����mE~V�z:˦�TR���ޢb@k�+eg���b�gVD�:C���`�ᨙaݪ�@�Q���(p�b�Q��t,�����	�x��`"�8����U�-`(�lט�
���Ėē���҇7���H�^��}������p=�ƙ)���t���ب"���.��E08��&�b0q�tð��|B ����rڡz6g��c3��n�����2�ݱPN,;V_)�[�4�,;�A���,�?\�Z���@|�>����1�~� �
B��5�6Czشj/�9���
�����FFɊ�3�y��0�
8_���]������X���l�?<4g���KK�[�	P����=Ӆ��p|���"�ގ9�4S�=���x��՞������� ��v�!(>󭁭(��j��河�-�_�Q�r ǚ{��#y<kN%>��#y]R�n����_�t=���$����U.+�U�#���8��Q�M��,o=_E�i��ќu�j��S񎏅Cvi'B�:Í^#�S�i�������������4�����[*"��ZE=�yf���_�[D�|��ɤ�` {�ϡ�@a2� �x��mF����
�o�kj��ʺM�k!ى�>��e�<?<�SFP���x3��y5;��s;9���Q�UO8�;i.�1���%���s'A���/�ht�H#�+��	��~vD��C4�캁qs�b=�kʞ�x{�������Z���[�]���qD����o3���@ǫ+�y�"������k����� �F}��;�.�i�uJF!��b�*�˜�岺pa�����m�E[�;��J� 7��1�<Y+�J��D�y��*&"F��G��ss���Ɩ��cO��P0���YB��x�����ؽ��B�\�3�����09o��P���s]���������������M��9�-,���lӉ8��΋�?-�ǹ�=b7ia�QJ�a�a��$X�^�X8ҝ�~���_�&��c5d�]�X����!i�Ak?]�2�[�]�ٰ��79N�RTd����C�z�f@U�h��E� ���`�:��<��B��O�x;��
��0wB9m�׀[����n�:Ŝt�l �_R���}�\N��v�x�]sYmVYU/u�,������?�[H4���oI�'�;=> t��\@EM\�٣Ӿão)V�6|%�r�fŮ#�G~a�e=ӃQ���4��$o�~l�Ձ���IF�.j@(��L#�׫Q��xQ�-)�(\:�q�!�g�++M�5���~H-69G�t��<��~�F|w^��2��"�M_Mz��uU:&��?9���a�������(�q�=÷�v붡E�xfa;<{��Yjr��# �:�%o���(��k7v�?���+��+�(+C2�@��%��kRh���}�B�ۜ����'�evObh�Z<��3�b���o�AS��U_��}T�9k6��ڊ�0����Гh�����h$�zՄ�n�^�ey-t�S)lBa���׽vt�����$�g��E�kW%f�Ea�D/�I��i����ů$>�lp��K���4�Иz�����GT�,����{�O��\܁6.E�t2�hD�E%'-%�O�E��!��u��l���s%k�Ћ[������ɓ�E)[��۝�-�/��	����-u�=��̈́8�Z�j{Q?���DA@�p�����}cº3*ʣ�M���*��6�-`����{V����Ś��R����lϧ���X�ۙn�~�m�n�\�.���.wB1�{@
����ÞU�S!Rh��O�a'<b=bK�8n�/އcnkߠ?�n����p��zHѶ}��U�L�:���b�U��9o�.�՟��E�(k�U	���^�r�TX<pHҩ���H�.�h��yϠ8A{��Y�:�9!k��:��R'��dO�����5V�[g{7���Ų�}�ٺ��.���ӟ/�@g:��w��h��9�; �����`°�ڂVx'=EK���̬�
�n.���۬�ҿ�IѺ:W�C|xG���|N!�4V�/�G���޿k�uVӏfk��dZ���u����˥�(�⤻�/6�]�e�ȄY�V:�l�N�q4�U^�j�#�oPa=�*����b�;9�ӫݣ�V�����&m�q�5TSc�w}�@��u|���%��wA()+��h��5���h,V��mj��]`'���%tpq��[C���A0�u��J)F�`,�b�'FEY��$%��(�oq����ճ����[>�qR���>��4�]~�+�.��,�|�}��J~��^�!�;S�5�_"�1�d�W�t�DJo���|��c���eZV�v��sP�(|�Vz�^�����0�
�]F�K�B��G��x�K�OJk�ݖ�ښ�m��Dp:��*Qc ���.��B��U����1�S�0�mۑ���x��Wu��v�x��fI2�.�5H�9��զ"�'3��$ ��0+�\�d:����N��4�1d��0���,ɭT)'C�I���%.мz���<�R���/������V�g%�'W��ٸ/Aܰ��i�SFk��L��o���[@l?ޮ����Ya.?|�$��Yn<���Lb�+��h�i!tjC��� +g�h����L�CX�5�NC�3�{_�Ջ�_T.f��n�aK0g4=l,�'֜-Zb��'��#W�<��J�k��83�� Ovv�nC�#�9����"��`�(����5�,�
ܱ���W�X#�?2oY�X�L�M���3��:1@+�9&�e�1�5;2Pg&����~w��g�(��N`���?�<��T��w�9ͥHY��ڌRDd5˟'TH逋�A2C�K������#ɚ��E�v g��������{0%]b@P�-���2�b0#��pu9Xo��Q�
��#�}���h��=�=i7��Yo&�!֗T��ꩋ-RH�L�)�����W��MBo���h�v7���b��b�a�R�^џ�oS˼i��r�[�_�O��b	_��"��(�g�@��e1Xi�$�`5Y#&���r=��]d@*+gF�z-�u�*o�8���o_~� ��j�t(����)"�3��]���	�	p(���]�p���.PsM�̏%��YI�_[���J~�m��q2��O��*b-3:�Ux���)��3�O�zN\%��j�(�fAS"Y�:ҙB�{��F�¡:摯�G_��BVG	����qP�R�����uBl��?�B�K���F��S�t^6D�`����-KB%ҠId�\��X�ʔ*�����AV�U�S�5�&��>��l%�ɥZ�9������� q�N�S����;�������^����ߜ��@�Bgn|�$ �tV&�Y�:JT���L5�I��͢�k���VDq''�EWg�ڳo�8�~b��-d� {K$~آHl�괭�!劼��A�G,�1��/Fm}�:��K�{��LI;�?�E�@�כ��E3��$��L�SM�LP���P+�RZ6E 6���*�#��5H�u�!�@�X�3.�<�_l�\xfCD�9�_��Kp&�$'��l<S{2�\��T6C6q;L�Mh�\U;R�y���sT��<�	�}�{�Ɖ�����>f�Y0:���i3�"
����0ýy[.E��U��Ze���|��ˬ
�x^땛J�={�����&�ք5ڈw�������@Ⱆj�%I�"&lA�����'}6��~�=Ni䪭ڱ�	��Z=I��E��^�;F���r"�M����BHc����C�-F����FA��i��#��~d�Җ�7pv�M�@D��&��i�/��Gi���ǧ������I�D�":e�
Xت�hf7���w�n�w�X<������h��,N��J�be�s���z�?���}6X���(o�My/>: ��D�W�Rz�*xkB�BP��/wBw%��%l6_�(�}�S]��YC͢�S��eVN~��5�5�c�!��-��*�l�^$B��B%&�0F�p�H)�rb��Ġۜ�:��$1��g�����Ǝ��q��Xl9����=�_����E]׎��D�������#s��
f�&�쌼E*������߆u�M�1R�LDA�PR��aP��3y�z{�ɘlE߹hq��.I�+@@��|3���)8���O���V�� Zoe!���LP�۬�>�/��I��
��d��B�N�����	���4W�U,s�-K�×��:�ܗO�������DYU��&&!'�*�I����t�\��kS"�R�L�t�Mu��*���d8{���ˀ4��] o���.��{����Dī7��e�f��n�-ɵ��Q\��� ��~(\�k&
@��mYȪ�D�ۧ���(&��[Gϖ[�<	Д2�iU?�*J�D3���Vn�o�H:��9��N�c�^O>= `�ȝ����&��#���:�=#�xr�޿*<.ge_��è��ܗ����f�p1gb�{�LpTF"d�"��%���N��Ls�\� lN�6��n"D��~���58��gs�q*��(y�Oj�V���%��0����uR�eR�&,���<��5��	
ė����In��w����G�p�r��(ӢDRJ�v?4�9�X*�'��ź��m�����->�[2D Zt�^�?F
 #�y%)NO�.�|{V�W�`��N�J�?oO�I�Wj��۵�5�P��d���F�u��<�Q�3fOxQ�I>e�Sm�H|þk���d�Ӯ}�`�H��ЃÇ+&Zc	n	�wn��ڏ_��*����שX�MA�ERs�'�f������!F 4�V�C �&�����:��_T�0U��6<Q�1��m�\�O暢a���o
u�t����M�nw��u�`Y���!�[�do��R�p_a�X��sF�`��C�����h�q�`@�U،�*�])}3�"S�^�Z��,��V�҄��פ��I�
���������ҭK�ء&`_����8H��q��M��N,�;yky���}��s���%���;qc�(a�pw�:`QmG7v���f\�?2��_@:G"J��v�\������i�
R��L�W� /[�����T1�T@���Nn�<e�r����r���S�t�����,�#�|�U����
�2�V<:.]Yx��ѷݔ��fSLu� ��#��*"��q-�@�>q�w@��9���؍,l��0Z�@ʩ�7s�@��F؋ !�joɸ�ϼM9�6�8�3a̼�-_���kc��6���Q��Y�;�ab�M��qi��H8{+�7���z��H�����ildS6]�aJ^��oU���7�u��EA���:S~���G����W^>E6��y���0��zN�ǐ����v!���"/��C��g�5���`maVp��=p��߀�D�q����@����p��s�U�_�Y0�I��aA��F.�Q�K���+m�&�KBL�qcئjh��쀮�,���; ��;I(����\�q8A:`��v���\;�t'A	�R�d�����������rOk���k�h
�/f��dQ��H�w��F
�eY���2YgCA���;�z͔i�p�j!�PJ��o[Pp�/�:�/�H;)iX�ʨ��ٕe]>\	C�	k��?!O�,%��1J��"�^5g���A
�-�54��30�K���d�{ZY'���AUT2�X57G�}LWv��$Y�(y����z��Y�x��w���ʾ⣤WQb�f~FT��>�\E��2P$�(ˑ�F9��Y⓯k,(5��<�+�m�@;Y�ZPo����Z>���\�B���V��3<��o��E� <
Y�%�W[��Z��ָP`})4@���L��[���7��i��a%��zu50��#�_�J��QD�$�9Aj��?z�_8���zßCX�����Ͼ	==u\�x�W'�4 �ƀ���� @;�&a�����1\_�	vg�M?I�j����Y`eo�"2>���Ff (���k�2���Mo�&�U���z���J����fx�����ܰ[	J���-g�c̫���w�%�
ܯ[�A�}��f�����FA���"a�d���V����� �ޠ�`]��nu��	�1I>��Oc�NT��e��D�m5FKg�^'�|��H#���QftҗV�ݢĹ4+٭�T�PPe�>��K��V�d��1��&��ɗ1����?�6#��qjZb����58��J�.�n�M"7u��Z����B���Mo쒷ȿ�xZoIao+B�,�(�����_� �{�����f����5��0�T�)��-a@YV��x���pO��Y(�!���h�BHX��������A�QN�<�Vф��u�@�dA^� �wu�fX�b��CC	��Ԛ�w>LI03~	a�z�����«�N[`�"�ː�ץ�4J�8ᛢ��F,#�C�D_��sH��q�.b�W�����7M��.�SFwV%Rj*V}��iy,��'�h��m��V.��m��jqo34��
U�lfj��~�G(+�N��(���5ЉG��A�9r �u�83���?�`���#���������<&�e[�4����� _�����6���#��$�8����u;�"Y���p�{DΆsY�����,�2���
�	�RNp%�#7�������?���ڈ�2��b�F�y~}�N��8��.�k�c.�Ӂ'����y>:��0��ht��v�X���A�t�]�lǺ�(]<|v��@���t�j�]�r���K�l��x�}P�"�A�O��;%�L��� w��|����ę�{S�f泚�I#���V����.����Ш!�&h}����scwmjS~xpl�>��� ���p[��RY�I���������bE�΀*Er^�1�!Q�܊�_`�O�M��_�5�!.�^�^��n�=Sa�[SdU�4�3o)�Ðr��TF,���#?'���-,@׿#6� �����O��A�v�iR�ģ_6:�ӁJM�}"6�������\ܔ���A��h�or��u`�i�4���(�uà�Z�=����-֯�b�k���s��|�
(M�l-Pl\��p(s��L�� b������p+�|�$(?z�LВiKқF`/NRq����X���p�4�^�	Ʌl� �Hx����TT�8�}za'#�]�+y<��Aɮ</���,,��iF�E��`�����`P�s�e���_���3m��x��uM�-�u�� ����2�q�B����#�G�7�cN�X�:���,{s&�Q#�S�큢�wHX�
e�蠁bz��rN�||�p�_-Q�Q�1�HjWK3,(�C�o$j��?(nWgX�����r��	����}Ĺq>����D�)#�>Y��C���������Mʈ��!$č]|�H38�I��b�@���4�������yc�:mL����2�^��"� *awW��B#Z?�o���s��b
��i�	T��q�
����awg�cti=�o�W*9U:>�9S/9?W�1gb��/R�h�f;;��?�b���#�Yfx�eڞ2�?��E&�]!s��N�9����F�Gwt�I1'��L-Q��ֶrk��<��~�@��+<�aճ�x�tg���^Q�R}�&�O�-�D�����hX�LK��V�\��}�[b#i.	���bG���%�k���ϝ*@2��h��gX�+�|8l����	�L�z�����LAqx�x�6f.>zqF̂�P(lm	��6�l�Ѿ��`Kfp7Z������ ���`��d1 �a����o ���M�u�3��|uS�j!؝!�	=��̧�V⿥������1䄲�$Qg����C��bM8FQ�2�l��}��j�1�5��~|�p��x��k��s7�JN�8�Ց��3=�ǳk�Є�&���N�D&t�ϐWS�3��*G�\�yܖ��s˗"�45F,�$�ղ
�3DaB��A ����]5D�������h)�}�t{�A�0��MAty<�Αld��&�z�nBhM��E�|�~��#�r#��F�c�Z` \�x'�U&.O�Ķ5��V���g���Kk�Ϣg�2���'�:%B�7If�H�^p̊�0B����Z�Z[���e�S3����H��Δ�p��ydAB�}�"v���Z5d�v����c�a~��WIJ;@�T����ζ�-�<~"�ѿ�S���u�!u:���R��(�jw4��@����v�
���es��@k�7��f�XA��
��͘��ī;5䵄��B���(X;W�g��Z�`f��=���Q��'\e)��/�O��a�(�RFk�+H��Lޞ�k���Ҟ/<sw1i��U�P&�Xbō��x���x��4���������g�P�\{$iR��,���K�;�n�&���Gu��`��BM���,طB+�E܁����V%�/{PE߰��3�M��9-{Yz��a�$����gU|�Ee�K /ڛu2�-��o�r�f��l�$ C��9U1tԭ)�lpR!*���B���\����Iw=X��:N��*��c�d�|��`��~]�߷;��g2�� ����Z��+���o�})��X�o|�P��ͳB�`>�6�p �沺$�<u��M8�4�h�`�`x��N-8Bp�g��=6Z@	pV<FZ,z(�k��/CP������ l�Q=*�3�~#��k�&Qǒ�@��+FB�M��]���%]M���~�&6�71���;>侤�22ǀ�����[^gW��وU.���݇�I|h6tn��"���ke�r�����]��:�w�cʄMB~�n��B~L��a���kX��1�z�e􀮤q���au�Ǜ��^�0eyuĨQ2���\Z�7l'V�}˜`&1TcJ}Kz��H�2�����x�j��]���߈�(
W���J����D���x��֤,b�Y��҅u���hBHL~��_�L=nA)�d�{�6��L��.9��dY=9��RBf��U�/��� ���5���H�x�`�h�4Y(��O���֌�o���A]5�ה!����B".dD!k3p�ކk�cR��Ț�6������&�]�F'��ݖ}��$˟[��YO����=�	#�z�P����kQ�u��w�d�Ǉ�k;B��`��t^�}�My���~���[���X��n"�+�cf�!n	\p�2�G�lUs��VG{p6l���M��?E��)����V��M
�U�x����.�Z:���z�#� g�_�ξ^��%�d������j�����5}��/M<QyY����6���8�1��.����i��r�6R�]9�܍07��r�7۸�����;r���H<w&����Ӎ ��U�2Ȑ��i�6R�������T)d��x���0�h��c+�l*_;�8��̊�1TOP?�~	��K%;�P�8���\�q�2�H#�*�km���J��*D���/N���+ƕ���1�����]�99^i��Hv,Ϲ-+��/��<eW7Pa;�۳fN�mm�p��k����̉��M(��M��OV�s�@��yf�t�M�.9�
MGmA%�ߘ��d�%��ܸ��^��]��HE�
Y�l�4�\����
g�ף%lٛy�P����S8rؾ6cÀ�#YGC7�M�����i]e��]�n�,SxJ�����ֽ��f ؓ���Gn[�)���$��4�ge�Wm�S���5��7�#�:����H$ �FK�áJ�z�.��"~�~��2���J�����BnX"���ոJto��Y�$����,7
��ͣ2��gR�gQ`{�<�U3U��a�/�%�N��ڮ��I[Ӵ��7cd�%�B��"9Oz1CdJ�xC4��({y������N,�8X�yS�+��DǮlz��|J"=�H��_2au��<��S/؃#��Lmm^U$ ��&/��Y���g������m쏴�����ʊ����_k��J�Ĝ/R~H��z�M�-�U�pZU��K pW^�-���m�?��g��|X�~�3�j��J���jz{عR*�*X�t�j5��%ͅ�ڗЋ?ۿO:4@�R��I"��]��,���G���x*/_ڛ$��p�f�!�1�53��˅�=�'�B�<e�.�i�s�n&��	��K���50��*��s>~�L�'����I���23ܞ��^69�vtħ��]��h%ɰ���h��WvJ8�ȯ��Z�;���U�_i�o��0�PUњ*� J�D���o�{.[K�0�r��*�joQƅ��\P���Id6#�T���UuZ�`d��q���FR�;��\S�5G5�?�m9Bi>?��Zc�z��~�TnP�×j������#�������MET��$R�������9��o������S�Ӧӻ�֖�e��X�J�~�C���p�������-\�.\ń��17���8ۡ��2b,���_�w��?H\*1�p�;_4a�?��M��& ��[	����*�����v;����7�?)���� �Y��M=���^�1�IE��Y�0 �w�H����2F�x���P �3�hDrb��;K����i�VEL��w8m��&������Mc��j��n[�A'�.	<���;�qn5��=}{��/G�H-�~��Cz������*w���;w��p��5��B��Y�ݦ�@`Y�K�������������p�M񗢸.'F���<�W���S��=+��/%�6��7%;�[�~�����,% "�'�U�����a�sL�"��,i�z�)�N�5H�)HQ��)*L��>��/����T%��h��)��Q��;�������+��H���UZ�D3�oM�Y��QOm��Yp)����A�����a��� 1W����W�޼��Ĥ�m_�&�q��.�x)�������f���Ns�z�W�����DKl��O��"?�'���Xy ��m���T��� TEAAv��7~i!	:������\���G�4��s�������^a���H�j�YW��c��w'Y���C�ŰN%��Sid�">q��qe�L��͛b���yg����4�L�R	 \�����p�o�w8��0a
�jz�Hl�6vwr���.̣���_@��1wC½����B�f���ܜ�dm-˿�j#��숲A�.��]d��yǎ������q�RB���,��PB��F� t,ɸ�;��oT��+�B�G��J)i-KD�3#r_8 ��1�:ͦ����@�c�-I:67
���^�-���*���(Q��9U̿|_���J��9����ԫ�A��qA�Bk��EAuWe�YE�27C��0r�9��Y���y�ʃz7��6��.��E����S�����=��f���b�ˎR��5�O�0�@9��SHF0h?�1&(B4e��������y���9��Z��a[ö	X��=����jP��M`E�u+��=h%�M ���1}�	������`��-o�oeu�����L"D
�������*6�h]��D�v)���I�c狜��=��lI�QNuJ"���va�4�8O�
��浂)�j����@T�L+�P�� � �d �k�lgG��s*y����8�v�SS�:���9�ę؎�Xr dB���:P��뱠8ʀv7�{f����q\�,��'�.Eq���\\Td�פ��"m�^�I�� ��k����A���cև���	7-�o�z1�|�-�z��s�[��t(B��;j	`u����@�krT�[�ӧ���L�*�2/g�i����,^�]�Xw��L����d�X�R�����4j�*���1��`M�c��oȶk]�8�hŪ&���æ�l:��0DknK���o�>z��߇��oχ#�na��b`\rZ7��u���E�k=���mcQ �-1��54 ��&���i4ue���#٩�H������U�?y�d�QL.zq_=��v�����˧BT�}�9��R<��gs29�C\#>�:'�8�9��	�}޲�,�/ko ��3E6L��=��Y�m~�7�K����#���s�0�:T7�k9L�X�,uՋj{��i��s�(Q�K��_��4�\ё&g%����]������Ҹ�Ɇ�w�M��*7�K^�g��H=?A�O{_�9DG�����\�V<���yeC�Նo3����R��#0���q�����? �F�B�(A�XL��2�J�8![��s$��`|�Î�75|���n��jo�T�fQ�s��bLL�Sׂ���>+��X\����sy�HvI5�Q/��4l��`#�i�{i/��Dw� D�Z͒�1w��Y�����m�Zg5��ނMN��S�ƈSy´7�_Xݐ<�y,�F�,�K3%m�E�؝���ͨ!�k�u�Y7�*�:�9#�!� O��l�����K3rc�J0 �`m�W=6��6-�����=�,�*sߖ���I<o�0;�Z���s�����U�Κ4�9*��#����%��1�����0�����w�m����/|��ak_�;�J����(�BjU��B�8�y���~������G �I����|� K����m!_�h�#n���O�[㭑�[d�7�^�L8���~��l �y
h�@�H��gY̕���눾˛ox�Fn�V�o�R��xY��q	d�@N��ExZ����`*0��.~#%]?kЙk� �C����#-��U
��>��m t�V=�\6Mb�N2"�O�B�B��M�h{*x�O���$%`�@cl��tq1���%|�����#֣G�uѓ˙W��W�>ʾ ��$H��/���Q�x��d���}	�r�rӎ'��L���@m�g�i��b�?1|�\�x�w��sK^,9�nu���3��M[66�5ٝIIZl,;��(�$���;�=��ɨ�1�^;��؃k�S[��0����~b�[d���4�MK�,ė��2���ɧ�4�6�r��tE )��W�׋���֦ �>2�����-��)N��D.�J�m�ʲ���e!���_)ݮ�O���ǂȅ�`v팥�z�<B�r�	1v9f��Aꡘr��OV?�]IB�2�Bݖӝ6�����F_wO���?41�����J��B��wLzJS�tN~�i��Ҵ;�Xn�^K�A(+\�\gb�FEk���O���]:�9;[&Ϛf��<���"��������L������B��5V�)���Ȥ�h�x̋ �0r*�2bЌ���m�Z��|��s�/:T� �+U��"٨�9�#K�41Ӷ�tF�o���.$�щ�ι�~��<0|`x�h$�Z��d�4��e�)����N�&��޲u&N�O$��BoT�B���� ��<h��@1����%��q�L:%_��qx��~���X�� ���|�e�S`�ӆ6@) _���1.�X1��+���� �����_�����mhŌȞ�\�0T��G��Y�=�k>Q��w�q�ߝ{oB����_^���]�#�� ��#R�EBw���7�H�"&j����
٤�RLϯMQ�%H�0��H�����e�>wpV���vgNѹJ[E뷉?�W;0��xÃ#�B�9}$�}�I7��.��X=�M�h|=S�׭D�W4u��]� ��R1\,L�ң?�t�3�R��x�'�E{!�����t�6/�i4��i2_i�Fcad�{،m���� �ǅ�E�� D��e�NI&%��E�hB�3N�Dvچr�,L^��+�YQq��!"��r��	m�E*D� �5�]n�zG��;h�f������A�P%�5o!~G�U u�&㰁텝���Sn��Ԑ�?̷��h���\j�v�˕�fsI��p�"R���AY�~�.^6>7�8C?p��:�����#'ﵑl�����o#�y'��)%D�y\�~��L��86�[j���Y��oFQ�w(�0" }5<���.أ��J�@�6�󵆐���X�A9�Ӗ�d}.��즌�?z��L�]��u  �u��1\\��A\-�W(s�]J�w���B��H�
V�u����vPfr]��wV���3�H�K�f�ŵ�ǟ���,C^V��%�;bڂ�.,#�)Սy'7��e�_��1�\��S�8Z5<"Ν�a�TH����`��I�@<.���07F�}��J��@c�zH�Z�j�{�df	�.�n^�t�w�9'��M��yF��@�~�/��f{��6�I�����Jk�)k}��)S�n���#�_kd��O���D��W*��3�}"#s���3�Mi������<�-
����o^�d�f���/?	�R�|����-�̨�1��u(R�}�G�����ϴ;��2��%b�y[0*�.�d�q&�T�F�1p}0*zI���m]Yt.�xy|8�7�LȺ�öC=��&r����,������<UJ�=<nK "��{�!��P�6��{����d$��+��d�H�q�Y���!��o�Wh��ݰ�2n��m`�Ѹ��|uɷA�[�&�X��$j+�!W��<Ϳ@�6��M(���L�N���1,e+��PЙ��!V���K�ΞM����q��:x��j�����"�KPv����xg9��{y�+<�'��m��U���;�xu?������R]%�C���G�Gߞ�Q�;�݋�:>���ڙ�eڎ�uA)���L�+���2�Ȼo'A�&& ��jPaE�K��L��n|-�q 	��b��1�m��6�&�)\3t&N�Z��)4���"z^C��Y�IHJ�}'g��1b�U9�-�,�/H
�0.�~�k�"�Ցx�v0�7�Sx|P�p3��o����>q[��4��^/� u��c���?IsX�jA���Iʪ)X�rA�҄��B��uV&��v��5!JՓ�s�}�.��|��p�/��V	���Ң��!@:���@�8����J@�r�?ғ�o@���<@W��)�W�PI:#X��iヶ�������!�o�����ׇn�#<x�,�V��48`�4ˇ�7�?*��
���Zo�)>�T�����(5*�L�H�~���CVJ��d����Ҍ�$�.LRy�,-���a&�Mͅ+�Ƞ�/�u��ܬ��<��p�guMm����}�T��1F�ͣS�%��J����]gA@���k�Қ\�.�V�T��Qm'H��5�ؽ%� �e�@`���Ǎ�5y�b�S��&���9�3��~>y�
<����O���.��������Ǘ�.+A)Ryä�
6mg2�Pc�͑ߘ�2�L���B�:�$ӧ8�KP1�]�V�������d ��ƈ9_�9�V��yo�R�@�Q��������5�B"&�.�?w7������>zV��۫U
�ܻ���s����A{��+��>�r�����i��ɱ>v�֪HX�x]4l�yLI���眬����:a�.���t�����'���4*L��l�aӧZ�L/�>w����Ý겐�\��t`cI�Y#�=ff��)�)��&��Kp�da0�{7ʒ����)Ʋ4B*�Ux[������5m�/�n��y�$"$��dm8�g�<kވ���K-K�HT��r���x�Z��7#/�=���
$�����)��S8�c4x�3x��L-kz].�&{��3��
����:N0�P�8�'b6����Bн\18���a�^=Q�6u�V�L��fݤO��xգ�3�O;�QQsA����|���������,kJ��W]8��O��0�HD�03N���@���XZ�;���L�d �(���H
	u���;a[�JW5��|�>h��wY�|L	�ޅen�݂dq��Py�ĹVp�D��.)��|�����JN���A=l�^yMU%�.��5y��Gq�h�z
`�!��x}^�Q�aZd^0��-�<Y�� �~�P��jot߰��1xWLHxN�8��2�qj�u�b����"��P���ỉ��`��Y��\��-T�>�WƎD��[`�ā�{_<ߊ�`P#��+�2�u��o�g^� 0�;a+�2�x��n�_ܐ����RD?�w�(��r?�
�e�̗)!�+�~�:�+���F̷TN��>x�ͽ)'�;k[$ ��X��2^�ȰlK����@�z��Q��PS&Z)���?i\Sqw�.�6�H	�!I&�m�����V�[C�$wb��UH��2T��X��+�;�ئ�-�M���o�X.�m�Ub �[iN�,;�� �oXv��d
�׋
al[
`r��@إ�=?f���{�<h6K��ec(�{�Mz[z`��{!]��$����q~����#Ϗ�c̸��=8|Q��uƥe�N�׊/p&]�P�3���pOn�����ӊFQ�����.�#��n�:!�C��d7P%�.g�����u�V�d�lA�wo�M��A7d�m�6,��X�'^dv��M3�j�@f�B q�~������ʥ�k)���V9l��Rԟ!΢���"�d�o���>Nb���Ƃ����V�|�^'���b.q�>����.�*_�D2?�(i,`B��%$�5�Ề�Vsdh���W�PG�cuF�L�,�H[� �����4'�kT��)>�u�}���R��z����}fk�*�ޜ9�}{7��	iqJ����^���x&��y5�_�m-qI̻��E2:��#�	[s,s�k��B�$}��%>p��v����WC�#�*�?�c��)ҔkV�A�.V���f�� ��4!	_� ��T_�=���\�����ty�53b�%*����ľ-�Е�BaM��{�eI*�^e�������"d֥F���&gX�g#jЪ.�z�B׹�@��Taj�W����1�bJ���"��q<���	�)�Z��Vf��!P�F�m��;�8�����vm1�V�~Q����i��nox�g��6�6�oˡ���w�J���H�Xc�|Zi�\���W{�A>p�@��:�*X'a�=�^�'(�͂�+3/B��Q_��_��2mKTX'�#��"��I�]P���p��%K�dd,�*2�F/(�뾯hk x5���w��<9����3J���˃j��r�ق�N^��k'1�{�W! Ȁ?ɗ�aS��H؇p��TmQ��:����bA[#6��K������uA[�loGI�*C$���ڕ����a:ۉ��@IP��} ���Mvs�i��E��n���X'�Y�o���S�c&U`m�����f\��ޛb�<}=��Y�|��HX�ܼ�J Z]������!d���i�겖_+����=?���:�F�PAE?MŒ�۷/k�+���Y�&Fq���(����מ4K���G�:���,�e�)��n��
J2V���[�'�2�}�*'!�*ȉ�����F��,KH�Gk@���}�^<|��D֘���I�'����A�^)�rh�*S�[��8+@��b�]:i֡*�O>��o�~����tO�R����w@+��
�bm;�1��6Ȍ�|pLp��0���������҅�Ɉ�r͉��^���)G)Kh�$�\�a�UJRru�pCs�jB�Ԗ32�����E&��s[�
�9��YT@��C�|`���;��8���Y�H��Փ� u�̶�8o&}:Խd����Y�q޾�U˘b�O����	�l6w�'~ֶ�rpW40�b(���s��<-b�jm5��)�N`��{ {ƌw�$���<Iuc3���%���o��WKiʘ{;=:�ZO[>��nˎ�>�|�/u	����֖0.m.�OaD��4��O�O�+t]�VV��;�8U��㴋
2��u�� �4���͹5������E���l�v��G�H�3K��+��V˞8��e�A���c���?����
,��5�&}P��t�`D�(�;n�߃?*��Ĥ	2��S!,]8�1�S!��dg	� �3f慣mh��v8����1G�(�N	:�e:G���@��� �dk@jpY�p����F�NN{/RqE�*��t�)�#�!�T��u���4��I���:��{�²���]��I3��EϏ��� �J�P�RȺk�V?؜v������C{���c`~^ht���`Y�Z����j�H�Ў7v�Ӄ�h��a�gR�1�6��Xy����y�j���u�1ExC�I�ύ:X���J�4)-\D���U���0'bi�q��>r$K +ez�d=s��je\!J�ٕ�~��z@L�;�\T��s��#��KG���O�x}06b�3p�2'�q�S,f�62U��KIs��'����g��t���^J$�p"H,��^��J�_RgBb�W �س������ώ�1�ul����CS٠(����"2!"B�z�Dޓ&P6Œ�N��>�PA�^хKI)�H3;����
d���_c�<G�I@��u����?��y��.�h�E=�Rā�2+O:�P������k$|Y��\��^�GmH?�r��I�$�Vvx�V���
��J�L�|����IgC��+� ̦���U��+���@ԯtg �ĥ>��`�f����P��˪��i��/:9��x�����#�f\�����U��k�}_nJ<0|���pSގ*25p`����B�,PF�b����<5������aa�'�$����)ЫxPd]�gQ��#\�Z��pR�1����&н_ӥ�o鱣CM��/�؛[�K�ܨ�1@�������!ݯ��O�|�R�ID��c%
�I�7����x�hL�KV�q�)N"�Y> =�����ϭ����ېb?v���ݺK�����-�X���>��`8T]�4.��:ȓB����E�\7�3�1Lq��޾��pc��#����ݬ#�B�����/��e4ۍ������G��D�FD��\&�\�:�a0�����"F1r{�Ջ{h{)�e�s����eV6�@����Źs��TĒGWi!6��S�<��a���Y��
�at��ݏ$�)�S�{b��M��������v��� ���"���e�~�Kψ^I��b���N���`�H='��Km�ϱ�l���do�i�������X|���אp/0�J�6̳��)�HM^�6��[Q��y�9!'���ЀyE�}zX�L����o��:���i=q�����ک����������\ *_X�N�Lv�p�(�4 �^�#{%�U���'��e��j�o6&Ź
��\4�y&�����2fS#����aP�S�}�hi�iVp���L��m\4���Ī��B/�奸�eb+>c���(N�Ў��Z�b<�`�~�GR���䍐(͌�l<xD��Ǎ��:�}`���M�ɒ�[\Vb��G�k��81W�$�j7<�|��9U�FO)J�$#E�u ��(b�_�8#��0�!;�*_��DZ�Dj+*kM�~�>O��#OG�1�<���[OjdL�X�T����u�7t��рܜw0������R��w� s9��>P�>R�i�`9m=]�&@Ϻ�#G�e��u^�s���0̲*IM$�T��f�=��I���uΠ�<f�v[�=�k�v���.L�Y��"�.�(��aL��l��Ni��
���07�z r��*`^��$�O�S)��4g�w�J��`b��@7:0���& �U| `������'7�ev�+�OسK�=(�5�.eʚ�`A�ǧ^�/�������������n�z ��D�1���S=�o/�.g�IاJrϮnD�cy��,W��NE
��НI���C�v��Zji姲���J���&Cb]�w��T�#F�01G�D��'��7��ZP��O���M����H��=��� WP���?�/4�(�mnS�����\�����)�(�:*$B������M��R�����v�xH!���ږ*T褡k'(�H�HT`��~d���:�WID��%��9H��~yj�놀��[UPͅ3Ҍ��,���	�3O�rQHs��I��	���onE��1���*�p��;�Q��ۧ�bV�����Bt;����|?����&FL�SN�'\�m���J�V��a��:�~j��/�T��2v,b�|��-��ŋ���
0~�fH�$�J�$x����De��������������?٬���Y�̖aИm���Q%��P.��DC�Ѷ�̦�&m�Gz�D���T�~�A����� ��]�n��t=�d�M�ƾ��I�v<��W*��u�赥ŧkw%̽�цp�}�y�-�c5��`�2�z� 
u��o�����R�<��xne�
Q�$OEr�K����hF�;r���ܓ��f��I�.0<��۶-q6�^�l�Ty�Wa�a�?4[������%�s:�U=�Z���Hu�N�� r(Y�W�=5�wG��NDMz5�w0ɾ_��_��v��ݺE�iXr�xD.U���tM$�^�m�$�Օ��Fk��j�o,��:P��ډ	�$���{����������w[Ғ�W���ED�a�M��C����(&��̻��Fa?��#���鷃kfb:Jg4�%��n�}R|�Ș��AY�/�e+Nl5*� �<��� 0w
�~n��հg�:.b��,W��v�]�M��bg�{�vogdK�s�/�$���2Ossl	U���#$�\���:%��|��婙ߑU7�2�
�:#F�����4_
)�+l/F8#�h?��%��_�!�� �6PǟN�`���΢��~ޓ/�Ϙ$�����|���ۦ��Ⱥ` }�s��]A$�|��C �ͪqK�B���5%v�`�#@\Í�f�hsx�9�QY$�h�1����w
���(-ö5�"�γ}�u�����E���AK��Z4�p��O�&������&>�x��4�"���=�=ϲ}���}���Ӳo�����Q��"��[{u�W�f&����\$���NX�	�����������y�:���>|G��T�2&9	��v�uY��s�Mzgف���a'ܲ���.~4������x薨ь�(���;��r*o�(��!�ŗ�@¨:��[�9��1wx�?��Q��ߣ�)0���ʀy�E�ZR�#ǃ�J��)�EK�a�uFl��� ��s<ߒ�M��":5�7KB�MT|Gx�qhȀ�6��&τ�r��K�Rʪ�Y�U�0���$��E\�E,�]�z!y�j���[?HC<�
Sۅ��h��s�[������=�|�fU��I��� )a"�����M���^���r���%�E�.<uf�z��?��^��2ℷ�߆���;l���7��1��=��.-:��l���q��*X����3	��l���c#l�(��ci�Kl�o��		��F�5��C��`|+Y<Ac�ab������Ay�y$Uu`%V�h��ط���/Î��/@5�/D2�$dƦy��)|.B�m���v�����i?�W�FX����ɱ�k��NlPo��}�
�J��}�ˤ�-���s��[ֽQ��N�$�������������4>}��!�3�D?[f� @�Y
��	�YN��rU�`b��R(�C�� ��F�-�H�u�ɺ��7&���[ny$�̈́w��|��F׻ƃ�m�f��������Ku�����&���3*�0�uS�$K�S,x�?�c	>�Γ'Iҭ�@��j�OҠgfA��MwD#;F���0������Ҁ��t��8��=]�l$ߤ8'�,�?�NЯ����������_��4��\3�o�ʜ�_�����	5s�`@��k�"�sS����g9�3�&��2`s�Z�c���r�ހ!�b�t���'GB N���|����vӥ��e���4;������g�*�>�5BQ�Tap(}��i_oqq÷��M�i�����1��+�.�^�o��\Tmt��sƽbi�Ri���L������N��U���{�fK4���	�n���uT9�n0VsE0&o�������0NQ�R�C�].�P7>ץӣv� �H�l~�B���a��{痝��$��v�����[cu�v��BD�8�_58�se<3,��;V�X4˾� �?#F��lu�X��H��z���TUh�e���l�F�3� �Lr���]aJ�mR!_�i �z���Q�VĀ�6�V�	��
-?��&Ys�/tw5��y�e�Ow�����:���Ņ�m��'��P�TH��{	�����bR�/,�gZ���p�2���	o�t�`�� mo�)qM.1q���<�L.�W�3�򺈉�K̏r|�a�,�?:���7c��q!%������]�A�<ik���d`�;4K��GY�,c8�H?��X��{h�K���^�bv�+0�aw�:���腐!b����";c�����t�{W�'%��
��~1MI�� �}�?bm�9�Z���_��'Ƃ˙��]�^��C��1f�[o���R�xP'��)k��@]������Z"�kK��Ap<����`_ݩ�M�L�����L��D즧�(!l~�C�27� ���������c��u�M�v��}���VO�*[��FԿ�4	Y�����&xD���Y��0��bZL(,�^����q-M]�,��:��@'O;�o_�Z��w-�����x��{(*@�7�SW$�����F�5�T��/Lt�σ�/vB<*�mx���LD<"���K!yLOJ��(�2t�*��*H�PN��g0Ķ5���Dm��m`b$�7��h��t�оXP��_߮z�e}���>8iQ��*�m���g�Q���N��7T�d.M�(��=n����Q���&�\�M�k�B"��}�3���g�0¶��H2b�O}��� �.���'Ҳ�xBU�bE-VR~��4/GZzzG9�o���0.�MQ8�>��yC�@ԛ:������aRF_��g6A��͚R����8|�m�ì`��֩g.!E��Nz$��$��+���/m^�t�dj��T2�͈��ӎ�����WÛ=��;�˭3�o])�K�x��XyF�����W<MWJ��\?ne*�?p���i�F�!m������f����>��$�$�;�u.��b�/E�L�&�)�lA:xt�c|�b�Tm-(�и4jȬD�q�k@,K���Ł�hU��(wY����/I��WD��H�4jP�mIPb�ڷ�����uAe��w۬/'B°�9�yO9��<܌Wu8���FmZ��ߞ��D���ezä���n�6)#S�-KzC=
,�F��Ru��c�/w�#N��i���V�RQ����"=	�KQ��(�� 1�Y2�b��hKH��7�!Ʃ���u��$��둺�b�˥ߵ�⑙���8��t$@�	㮜A-i)�"�'��٬a�4�h̒��W���T�4�`���[Wg�t���4|r9E:���S>�DX���ɢ	P�
�_6�?���@P��]Y,�vRYSoUQSH�KF�!���ҩ����Z��O-�� �<���K�n���2���]5$�+�/��/^���	�]�bNۋ������HY��(�怼�_'��'���fZ��QS�;��4�8Q\0�������3{����}�ā�a]�Vl�k��j*���Jq�i M}��GzV�p�5-�E�x3�90**i�W�o%�1-��u��K��g�"�Ǽ(���V�VO,D4�	����nK`�h��/���'&��6*�w�j�:�RDŕ��Y�/c�s����~*`��(���:\�W���_��'l��b���'K�v� �& Bx/P���.�U��;䃅��C�Hm�/��}~5K���٤ �w�p�j�ڎhB��i������:!��TG��e�Ak�Փ��`�s�Sͮ[�|��_o���N<�r��Aa�9<���u�p��m�'�I��8�l�!�eH��(���k�y1�a��F
iX��I�t�05)��=1��e���h��������VP]��s�]���Y�c�f૾�}��hj���]=�åqр2e�Q^���z��ah!������3�f�\FH.����Զv�#�L[�l���u�(9��9�����E�����G�D���ˤ�v��i
l�l��}q#�/��� nVD�Q�F��MS^����٨b����������k���g3=��QR�iY���@�0;A>���eգHy5O��
<���B<��쪚��&��(����3R���z����������]G:�}�	XK��:�YI�[0�B���XK�J֒W�֩ժjLY�[Dr�c�aAMjɢ��&2;�Y	�{�3���Na뤎�8�,��1L���A~���W����feds��_�3_b��Y�!b+�b�O�7���s|��۔}�'W؅�g�uLD<;���wȌ97e��f�� O�!����7�$t�u\��������x�E���:f�����ۆ؄QFX�	�yRxV���Ax[�yj���RZ��k��KTg��"~�㡃�sT��_u8�L9\t_&���شR�~��Kz���q��H�}�%U�-0�1���j��_�GY'k��O���#��8cp����� ����t9팾���;�&ӵE%�\J������W  ���aː}��`׽ۤAѬddr:���.���/�����PKXlf�a@��V`D�^"˳(iY�R�:�i+R�B������;�缴g�c��I �b����o�>?C<
�z���h3V�G�%cj�[3�ӓW��^3Z9�|�7ItZ�C.ǥ ���ލ�W*�%��0yTnAW�I�x��"�ѭ!@9��h��I�4�ag���G�hPDꟍ�s��n�w(a�H�צ����*59Xh%u7m�+��_�dm�VК�sZ ��*ݰ>�KI�?o"�P���8�\�P��>7�2����z!:Ƨ��k�.�$���_�w�T�'$2�K��<Z���3k�E2}Y�@��α�$�D��մ�B�j̚j���8G��h�HdF�'E�G~H��m��T�ܣZ�ai��_�Z#b��� �ADO���FS�u�CA��|z3�G0���.q�(�ܬj�����WlJ���Q�1/b*?���ݤ� #V�ͶP�Qg�m|ԧ+��c���!��=Q8م��o�YsN��E*y��9�"�x�D����e
޳��)�d/��0K6�_�>#�B�1�|�g��*�%D)�c�7�ٟ̚�f�x?�߆�ˉ܊�D�mvd�iA�cH_��A�H��0v�y�8� ��2,N$C#�;�|����W����`Hh�{��3�F��r5��e?���D(��<��֢0�./��`��|�'��ᐓ��[ms�[Ia�hn�s�0���Qu����G4T�w�X�Վ�.ex�!i��Խ��N��M�:@u\���m\f��+�+B
$p-�kSAK(ĚӒ�;��<`},z[�y������0<��Rb�<��䖁EUr��~�ƨ��z��odf����x�	�!��}�G_TI�7�{�<���c��	��]�%�Z���Q5&���&�Y���v>y�4���?��Ak=痲LJ��"kj�:�F/��0���
�)\h�}];<WP��z�)8�&r��q\��jt��~ߑ��.����Yx��/�#)<G$��%�M[��i��i�E �,M�%|�1c��T��i�A� )������(f��!X��S��&��6����IES��#�E�wV���<SVg�4x�=�G���ާ��Ƚ3����[i4�O�ţ�i�=�!��ݠmV� y�Q����O�`:��D�+�`@�����s��r��@�=�sy^��}�l�<���t\x�55հ8��B���`F_�Rv-�Mq־?�����������}�(�?D�k+_D�t#7ۻBE2���"����{��^v>&%� NQ&ި�*�Q>3O�k��P᭓
 D���;G��@�ڊA[t�VI�����r�}61g�`!�=�|7Q����kS�
���m8��Ǒ��ĘA4���hy�n-�\XL9<�t,7�3W*XA����,+��Y����ᒆ��z{'B�~q\*6��dY�R ���>��5�Ż��ܿIx�>�-��>e���)R���_?�u�YZ:!R~*�a��X૫2D4�n���4�_E��/u���]u��6ؖ���gߣ"V�=��Aǟ�iTv�|5<bc����R'?�∇Ҥ:c��?�Y���Z��w%�^y4��6a���S����"�dڗ�O�b׾�7&7���
���<Й���j}ɰ��K.�!�v�F�&\�y"36`f�8Ϩ���y�r�M"ťjS�)�5��G�����?��,CKPȰ�h�b����u�D���:I���$��3J�n�^<a+M�!&:���{�&ힺVYYMVH���Y$�C@yX����¨;@c[�������\oI��M�F�UhZ_��>B
	��i.�JE�pi�2�؉������)�]<��3���\�sp��XX���)�/	�-@Џ�*�].�a��ڕ?�q�ع*��Y"ȸ�q����~� ���A~^��㟉�N|��}���ɕy$�a�@�3i����@����Z6� EE^�c���I�Cn�:[��7�w��P��-��m���I�\H&̐��h��-��C�D��%�
sIq��ڰ�2w��{k䉨 �_���G� �/�SCJ��9���+������m~�,��]+v�A�p��r"������1\��M�DEA�*30;/�~��B�\�,n������׫���~nv��$6$}t!����~
���8�c��lD�ʃk#T2J��a^��T��l.Ӣ�Ẍ́E�u{�ȍ�=��e»�K�A2K�Om��>V
~-�5�(�2}�H����H�1�W(>FS9Z�=��G_+5W����|�A��
�f7o��|L�t�:v�}���-%�FZcF�4Or;e���ֲ+ �MxJ��w%¸T�XG�~�zW~�]�����|\�'��5H�b��{���!E1��>�g�y۔'���ъ"�jy*����7f}����+��]ʭ����Y`�aXq*40�켌G���V����p�eU�j���,�W^���#�,H��p�߹&����ɓ�jb~�J��Y��2�eB�(��"b��[�RG��m?`��nKs����Z��_���.��nD�#��M���5_��q�J�c�Eܿ�������x4�����n�"�U��ʌ�#�`�)���H��X�g�X�沱�Scv�Ow�E3�o4ɸ}E!ǹ�.���[�����/��D�5@����/�mC��A	��L�������
:H���	�gh�xpO�'�]���i�~E�XJw����X^�0��ٞ��#�*�T3�.�×���~5���D����	��5�}�\����C���=)�ո���Z���S ş�!і��&���=ܦ�Ѹ�{�B���/! 8A���^.=*����!K���X��j�捚a7��@�A<q�tH��%]��MbQ��Q�O���n������p�<�s�c8�1�>��C�)�­��
�TZ�b"��;i�/�G��B����F�֜r&�L
	�į-��	�瑌�R)��|�uX��c#\�{��ۘ�|N���iU-�QX��DiN;?���'�з`�P\�U�E��+�V:�Y2Z��Rc֕G'  �;��� �;'��=\A,���r��x�g�{8��d�m�q��蹑6X_��$&i9-��fQel���O�͈M<w��%���_�|��H�Ȫ6怚^E�F�^r��^�V�Cԛe0X�!ʞΙ^�
_.���I�N�<��Gļ��Y�Ŭ�Y��������k��╡��F-��&�P��Ї��E�t��G���S�����K��� 	��e�}�0��O*=s��Zk�U��?Z�fT�M���+~c��'Q�Z8Ns�Y�k��s_?�q�f2"�}	��%�H ��9�
�LI)jas�2�:�X鼧UF����t�Ż�����JO~�LZy�Jc��[��q�k�W\H>d�bHO��~����ZJAK]z͐Ra�1��RR�*��	�@�M�/�-�~�14�;�����D�p�8�idsͣ�]��>,����}?�������r>���� q��I+ׯZOS�y:�ђ�?��n��x,�j��ހd�.���������W�� �%�\T�:��̙�����,�Y_�w�pl�\�1��'=L�c�$���!��"N���z�A�=�6���?�mԣe�&�I�%H�N���ЙLԤ��
@��!5�7mؙ�=I�O�e	h%j�1���Le� a���0��1�@t��)�f�EpM�ȝ6LN�Q�7ߔ��%K�V�\���Hit� ��rV��7#`���Ix�.o 7ۂą����|7�v~ׁ�D�+}@�S%��n}�݊�?�%���T�*��w+������U$k�9�?��Ǽ*�Z�:�c���O��R�Ún�����~�]ꂣ���f[�{:��*X�Sk$�.�o65��<h��AϜ		�nҹ�Uf-��7״{lJ�.'G������.�N;K~ eU#<s9U֚tfhf1��@XY���X�{��ɒ��U�T�0��^a���¹ra�C+��k�k��L,魳*
�9��p+
�ٿc�:�^��n��k[& �� �R�����y�:�(�h�Zh�!ظ�.��jr}�H�]
����V|A�z��g�	�~�4��}V�N�VC&E������ˀf���D$9��|�9rP����ؒ�^�sN�Z�K˅���C�pԾ����NȰ=d+��d��(F8@�#�hp��"�	�p���;���|��UncR�-#0>��c�(尟̻�2�Z*M�bK������ʍf.�2/��uO3�4��>�w���=���G{����������J�㬔%�' #�����O6�=�M��1�a0t�j>���*�UN��'����W�%�K�*m*r��p�m��Z����wo�[@�o�Yi�s�?�@|��\oeq�쉳؜t(�~ս�$e\R�]>�f�b��j�"��6aE�����B�I ��G�h~H�?j���I��i��a�9�����A��G�����S�q$foȠ�-Wlv	�qlU�gl�[z7<�w�>��?��l"4y�..��G�{�"��WI�I�W+�ռv�S���� ��g��B�����r�ے��2'�����;s�����	�y�*�-��5����F*U@���8�V��;kז�V���8s��s�q����2s��D�`�A� �!Ǽx��,����\���I�C�ۘ���W�VJ7��!;������=���\��@�Vfo;Tk������Q¥�* ��P�8�w�+f���o��U�Q�ur��ؾ5�@�0<ƋA�\��:~��;۝۹�{֒�῁��h��!��������GƏ���cA^�D�_d��	P#|�}��ǀ��,5���!�Ł��6���S���k��I>����Dz�j���w�	:��7��K��]�S��^��ݺO!�\)��C�I���}�0����	�s4j�ZZ.dMVd�l�T�xn���sAޗ�v�\��b����i����yj4)��s�.Σ���7�H�A1d|0���2+C��7��8�<,I(1���]vI�y�~��Ýyŕf3�H�c�ؔ�DOQ�{�J҅ro�`ɭ���	���'���H(��8��ʧ�����%kaOF5�4��z�(�l/��~{���xN���V #{��6��F���UNQa�'����a'[!]�e�(�Z�~�ay���E��r���j��S�׸�z�e�����H�b]O�ޡ�sɧ���0�xa�.��^���u:�`+a�7����ʹ[�qGP�Fww?Wt�w���4<u[��|�ma�2|D:�sOR���r���]����c���y%�ӑJ� �_+��}��7�r�%=�q��a�@O&T���S�vi�ӎ�r+�v�ݢ��-�)�Y��,  ��Nj���J��M�ì��W� �K�~8O�K�j$�-�anޯ�^�/��%� f�!sH1���ȑ5TY�K�8�Y���*x[i�2J.� �t�� "�P�� 7�b)��`L2X�u����b�T�z4�*E�h�]�<�	yT�Iu�z��;5�������z�"���z/Y���,�?�0liy�)�V����HV��]Ȗ�Y�[�C�6�D"q���y����ԝ}x���c��Wo	�$aZO�$�M�:�g#5�$�\Oy���0h�_uzEO8�6�`���/�q�p;9,�K��L|Ё;BSZlZ��4�ez��M�y�S��'s�Η7i�8Z@"�u������+>�ͅ���]����q�v��)�k*� ��y2�t���r��g�Rn4�ᇫ�j-��.��q��h�Y.����=��r� ������{NH��1��@�02ڻ��ށ��9��wH�,G�ۄ�yOo�������:�M�����_�����ƕ�'��5�#/w���1���jrSX��&��;���AM��M7�*��8�#��Z��!*M�<������"�k�>Ӧ8~���/(x(̑*����,���{_����*pfcy	�H�T6���ՔD��u���21�c?:��D5	������̏��+��y4py?U�"�3B������&�� .+n��9�:�^�	������Gx� �Fq9K.���Ȳl�����~�f-}�_m����zQ�"��"`ʊb.O�%�Yȿ	I	Q0�,�Fh��B?�T�;�õp�ه��0����s�����R���/x��!(�&��)za׈��<��O���u!���W�&L���-��a$��6ɝfD���D���S��M����`4�4}��'U�8N�3%�e����qG}o�5��PY"mB��AΌ8f-}'�A����ҝf�B�O�����@l
�	�k(�6,iXTǵ:1P�M%�����s�BB�^N��H1�y� s/��
�?|;S~�R�>_�/C��	g%���N�H�DD�L�B��ӊ�(Sg\��e©��z����K��^�k��U�=�A�V�尭��$��*r��o�_]rĲ�|���1r�����2�˷��{�8E$!2B��}��`c�>x��.:�x|�A���7]� D�<���)_QDΰ*7�L���M��{J�tx��K�[�(l�h(�t�lᯀ���@6��1�5��H����X�/yT	t�^�Rm��We���?�-�:y}���+J̵noD��և�)ң��~l�5]�©����:3�R���w�ٻ�Zp8�����OQR&��{�1f��%'�t'�l���h��E�������Ca�Ha����$r&}ü��v���'>������*9[�ѯ�
b��$��>1��+����!w��A��ϱSMo��7��8m��oﶿI��\c���R��l����9�2#A�Y:�*����-�Oq���U�z�в�d�8\�~�w��] ��&_�>o`�"o%�=��$7�����2+�q�~��s�.5�6�3��y�����g��]o���d�E�Lw�j���j�����K,Ł��Tgp?ߛY	����-���5�y�o�"_�iT��Pw��ldPS�A(���l�T�o����q����tV6yt��|�⇗kķ�ƭ�/C#4�3��3��+������ �$�Ϟ�����y��v�	,69�����ly�-�J=OB��).�A�ce.�,|^Tݢ���8��)S)\vh�d�*5ע�!(���{�e����"r�k����Q�b1�X�ר��}9���i��;��s+���8�0#�V8aq|�-�6\�W��C�GM��/�ѳ/�"v�i� 0���^���X����rѴ��rqY�o���c���"u55�+1?B�B���WQ�$����_=���Z^X5�h7�k��p��� 
����	�o[���A��x �/��I3�9+p��1���W> ���e�K,H#�
�.W.pd�1C,�۸�Ϩ�8
)�ݪ��~��ET����zԫp|@��AW)y�W6.#�o,yJ��X˴B���=���t߯�%�s�>㱹�\�Ջ]ۦ�J�}@�.b>���᭜�b|����V:

�U9��_��|��'֍�a�B�d�v-�,������(��e��s	ɽ;t�]W��O-��y4�Ѷ����7����`�!PA�B(�\�n&Y.$�G)�d�/����w�Y0�s,m�'��k
��V+��*��:�����B� �{=�
/G�;��~��������8�O��!	��J-0_MO	���k۩j逴
�j���?]" c�B�6��^@+�>
�}-����c����`�*�OD8��a���cQ�����׶J��ln:�t(��"&�/���E�:���f�K���d)��/:&��:*�.�]Զ�Rv����)���	��B��K�<�cn ���CJu�6��v_a����K�/:Z߇/*�z'����I�V}�M����������|R�IC��f��.&w�<T����%�P��o-��}���1�����tR� hNM�b.��T� ���1�%I�C>:�0��⦟�����T��?�TK96��y�l��6���(�&8u��{	��J��yCU���p#2�G�;WOԁj��p?�h�R�����T������9���£$vu����!Ek$U<3Xg������Tj�aJv^)+�ˁܵ}���w�lx��[z�+���t�?��p�d��WB5��������y�y�n�P��
4x��)/���������5<��+H�D�e�>�7�L��,R�5^{�j3��R9����a0�{�0Y� 'ʜ��~勠��RA�ޟ�Ma��H頾36 �C�c0�~�tl��:�G��S:�K�J#�&�����wG_ӒN�<1=%`!��OMΆ����$x@�����2t���.k�Q����w�_�t�V�Qʽ_;�nO���0X�����z���Y+���<T��� ��>>�9]���Ŧ�����o2�X�]~���Q=!��K΃kۙq�����|/e�m]�G�#��]k����;D��8��:��%�����*�A��/5Xr�p�
��_Q<���"�� $P��Ȧe-"�FI������f���4����uGǱx��#�k@P�0��"r$����u�K AF;��/�-�e���ؠ,�gnPZ�UH��/���,���[��)a���`#�?M��5��-G���
�@��YW��K�g>�Z�*ߘ�A��2"�\H�@ol���N��q6��b�UE��ܝA����DT���G��ݫw��Gd����Nr#�a)���|���z��@Ҭ-�7�]�E������[��� �=j-��'�s1ތO���RWK�E���C[���9���ć�_������4�*A/�<��k��X�o��F۪�vɽ��[�7����t&�03�f�9'����\�ƲfW�o`bzK\l���
�?�%f 1�ډ�bT)�KO)��1Q�T�!�3���˛��G�f��������7M� 8׊�>ۃʀ�z�R�TL'�� Z� ���fH�G!�'�Q.(�c���o�̯�)�=S*�͏�U���+O�`YM� ���2�گ��J\;^-C��p�E��xە����e�A:TLi�G~�'�!t�e�~��GNCT|rE�޽�"?�O����)-)���4a_����>�kQfϯgTܹ����c�B�+�M��x����Pw�S�g�m]q�������#�a-�}���?e?����j2]G�K���ٴt%�V��]�L�4ăi�-�S'z.�U;9]F���f��.����Y�0aǅ(�k���)��Vu��d��s�Z\���.��vy���);��#�W�/v�/�$	TcL��a�V�39.�`����aBVo,P��;���5�m��ڈ����N����Kt���h�m�w$?cב�����rb�5�mI�����L���"'lCe-�J��ɹ���^o��}}C}7>���� <��b�=ɜ��q��^��[���)�B�e9� ��d5>V1��,׶��ņ-����[�.X�'0����%e����`"�r�7M�8"�	��-ӸZ�,k��-�I�G�{r�f�i���)|�{�T;�[u^���HzwE�@�;���#�`Щ��Ř��]�}��&B�OC���j���	[�-��R��E��'a%�-�H���c��o;����~��	�8� �J��T�V@?prsfR2�z�c���AeBD~S�ȈBeՆ���Ygk��+��ᝢ�Nx]�n{���P5�2o�,ڢ(2�&w�-����=h����m���-нJd���D@��� ?���p=�l��l���\�6�vW"�#�Ox�j,tohlsL�{3F&�����V�1��ۊ�S���ǫLR?s�� �ޞVt���v�B�-�X���~�����b*Jzz+?V�������(��'����_�M��D�	�K6���mPZ�A/h��d�&��3��?Q���K�|v`u�M�a�yj��2�ʡ����u��1��G����B�7�(i<M��=��p��*�>���j���+r����=��7L�N�������[|-�"�qh3o>�@�R���_�XA�7�Ð������[V1�c����{�
��S�I60�� �����1:;^�H�G?]#\�\ō�M ����(h��+��t�$NdV���G)�.�u�M�k������������~I�r�<W��F&UDYd?��?����	$�u4�����w6�O�ZEӃ�[a�Ld�5(@Ó������.��uP�����ů�J�4�DC����"��[�稼�W�T�1=�n�5�i5rx�1/	� <`�[@`��~6�]V��󗵁�j�x(r|lH���N�q�1�	��J��VK3���aV)^�~3v��;�A���`l�*�o	�V����x�x2�7�#85?_@L�'uS/Cݨ�����y����Ҫe,�o}�S�n��Nl�������aC,�bFJ���-Z��m��ʆ�K��1Uy����Ar���&��g�޸An����� y!S6%����g���v���½B��&<��������#xRv$Y X-@��m
���F����\��]ϛ�۠#�H�kؽr}p!襜���:��24��G����,�O}���T�6rC�^�A!��X�����h��k�VAp[��"
d�oR��>y�i��>k_�<0E`G^�vn�s8���Ng~�Q�O�%3��y�Q�WT8�h���xn3�*XZ����"��ݙ5��%3y4��ד�룙<A�B��|3Jj�u�{��f��Z��I�L��ʓ~p���{��G��= �6	��xmg,_��F�
K+�˱�	vوt\��֢ �����0�Ɗ>��I�LA���21L�j7��'�2	$BxS�삣���@ш+w��<�_IQo����xf�|����v#���i��*��*��^�����}�����K��o�=�Q�t��l�F�'zh��x���w���*@�?�@~�������\P$���d�3�D�����t���S�]N�G������4:���K�X���͝>6x6��ɌF�S�.��"���Ͽӱ*�����l���|�ƉE�C�'��)nQ�����`�@�%��.��S@�'JL�<���]��'xl�N?�}����;F� p�?�*��䅢t��;3�F9�Q�Kh��� B{%�JH��{��!l �Ss�p�y;�ʋ*4^ôB�
�漴�sLT�Q���o�j.Xn�MÄ��!y�'|��Pg��[�I[�h�AP��a#t��/�b:�9�>�%or�졧a:Qˮ���-����f���I��,z9K���15_Hٓ��M�$k��Y8�����+W����2RT�5п���L^� 7������B'	��������pb�,��'�o�^)���m�c�E�>�����T��5�X��X����̈=
pU�|���~ᶴ/؆q�-�_�p�Vg��'hlF�d�Fp�w[�9��� �Ws݃��u_9��0��H������L��<�x|�cBP��%n����zTN�?��\B��t�V��?7���-�ܳǤz �Ǧ����}_��_�k\c!���
mr&��cl�ђޘ�ϴ~��A�^))_��xi/���#L�1.Lג�D<%�,��V������ ���K��/v4�}q� ��:�j��6I;��w]�����B�^��ΚJk�f*?�5�:D�ed^K�&�����Na�1��H��Kb&XDAPu��A���Ȯ�:DF�o_$��~n0p��?���u�E�n�pjZ\e�.&��6u������4��d#2���,������߫����#_�����@��Ar�%J}t��]�(�-�v�`�#�To,K�I����p1����QA��*�n*�+듬�<
�o�ü n�/���RX��آy˻m�mFPՈ+�L`�.}cq�,3�q�ĉH~W�,���d�V\nv(��Y~.i.6�]�ۍ�]��Q�[!هZ�.��$<S,+���̃Q�V6t�|��x��h�֢�C��,���
����3�+�kk6r���a��1h0�R��Q+"��R����2��֞��v�0�Dd��H��,�I��Rk��މ��a�c���h�]�!C��Ve��N��C9�ŨG4D�x<�ml���4��1�pF<�M�L�&�ָ_[щZ�F�'��xG�Js�C7��5�"j�u����
9&UnT�����u�
r;�]^i41���i�'U���8<(���i���{h���n�.vyY����/�揧��$�/�f�i�9������p�]疡SLxT�<�8ND;��6.$f�>uw����O�' icr&yc��翓=-뜖�`gy$F��5E��o/��)�@M9Hk(ȕI����e��D��(t�?�:2�!��N����v��\�D��f"'��	s l�ۂPy��
�y��ϔ��x�Tl?��?%
~Չ~��-+�~�!{��P�+���JzS�
S���td {t	�~������*�F��*%G�3'���b+;���P��H%�f]�s�7��O���p�����R<GQ
đ�&�P�����@R�q{�C�/�	9�MP�x�y9��4�\�)��c@��菅4� H?ex{��j�| 2B�պ�D���&}�gLp�<�\��e�����@{�P��e�ّ��^�b����3r���E�q��(<�_�K2*�u
;�J��)�U|��v�����26����K���`�i(�%GMq��A���P]�P��تaȓB�X�Ĺ�
Ѐ�Ɠ�����i3\e$
@s�}p���`��_��`UN����#Mt��d�+p�-V��l��o�_��6���Q誤�!qc�/�+�0������KV��3%iZ%�{���L8�e[ q�\���iP�M�A�v5�A6�C��>%q#����b�",tO�
,���x�DU��ݩ� a���H���힨��k�.%�����t1ԯг<6��&��P�'u�)�µ���Ј�<�o��l&w.����@`�N���|���ѹ��S�3�^�?��7.���`���Bf��/}�@�R!e���f���쌖���RΊ`�=�CR٩�a�lp�+�C�A1ם�jU�����)��C/�=�
���'�gB\���
J�o�}�o�t�~
�M����(R$��A���5�n/��O�Ė;�V3!pK�c�0�z�}���m���ڐ�b�"%�}u�-A"cZ���'A�m+����<|�<A�ϩv'���&� ������p��i�{�nD����9'�zpA\�����2��S��}(ÿPYv}Lzl��]{��L�t}���C��"E�����	�k���E�o��e�.�@��s�pT�'n3��8Ln:9����h�o<�fUj7N�Q��+�����BP�1�W��+)>�b��Mb�#dFþ�O��4��;n-Ⱚ���@�`C7O-�3��VC#{g�����e���,�Gϔ-�,�3V�}��1�L"�d �O���oz�������JA����e��j�s~U9�'j",:c6<?w���ߌ�S���C���┝.�WF�ܶB����|-&����s`(���T�ԻOZ�ljJ>� f�����������3��d"��N~�IR+S.$
{��Q���r;�
�F���3�t?�#�5��h���y��(�d!:n�9S�B:�D��d7�j!�F5�G��#�5�5����Jy��k��5Z/���8g�dt�C�hB��hͫ�|�hΔ�D�v���g&�!��~���i��֓�°Nk�?Qd�Z1��*��j�i��z��j��T	�Il���P�CYY�H�6Vp��v�������Q��"]gxqX�Qd��8��kh�����&)�;0@�T�wp�"'JFAe�9�˜��aa�?u��Hlw�7�I���*	����S(���/�h]�F�r��G.���}��wI�fޭS�h ʄ�*���l[�����)z�T�4���c�W����݁�?�K`R���=�w�o	D|F`}N�.^�ɗI�U��f�6��ɫ\���ݛ��;��|����MB[����W<[��^�PLw��M�1?�xzǮ%�?c�1���1����c�|���	�����C�LUz�LN�M�'��������\�f������vd���:��À��]��
7�#|lXUUJ~!I�`.����`/�|Nߡ�O�$�˜�>�f�?A۰�x���PHsݤ5ëɄ7ý�WI�rj�8>�d��;w��}G9.��ܛ$��@��9�m�S���˿r^�+5^W�=hC$v2;��� F�\���#Z"at֢h�b�[��2��7���oim�mR�?3-��,|��?�.�an�Uwli�g)�xX2F��������]Ņ�`�O��(���bD��9��&��|�
�$�zC?1��M�{t�AW%-��,�����^�J���F�:�]��$�]�b�|�p?ZO�c;���10�-����-�T�r��zY� t���u8��>��Ǌ�g���{�?l���̸X�ht�]k���FQ��BeY���>��c.U,M aݣ�(�c��#�S�Ӽ2��5��Q��o�[� ��`�dZ<�=�(�\�����<u�&���
��6��2��k��7O�i�d�ث$��_���Q���%|���m4��W���p�6�F3^�M���-yN�� ��ׇ,�����6��9tD?��|k�5�;��4I,�G,v��s(kJK��{�-���תh3h�O���(p�Kn�EK<����q]��8�'��a�&�?��a��#�H	�y�3�5Md��*�����^}$�ν�k^Q$|�f0�ħ弳�`*}))kmy�æ�a�&��jJ��o�x.s�EM �V$	
�<J|E�7ɓ��f!b�/�1C$E~�����\�붸y��N<���].i3�z����w:�qN �
o������r2���T��Yh�]'������Z}�?�"�ؑ=-8J�{&HT�2�g�M��_ZkN�vcH��-77ұ5+'� r�|]��HS/��Q��r5�qz�I�����!�Tx_t�G�O�;1e��i�z�'��ap����|]�=9B��W��2s���:�r������W
$�PM�*d_^�c�M�}/���,��P�q1�^�oY#�ȇ�]�����L�XW[��F����R�%��M�^���<4�E�]��Dc��F'01D�k����.SG�$���0�U+��j��Ϋz�|@��T�\n�dT�NT�C�P���A��~%2O�����<<�u���t����u�ٛ���dd+��(~s!���a��$+&AtY�u�{	��mxە�9*
ۊ�_�2��;BW�*q��h{��}Σ�;P��6���#ϔ�]��L��LtA��
X6��M�|ID��3^ Ϋ�+��yy����`���֠7���\8�eS;�}f?Sf�����]�8��&��]�<��P��'i7.i��.��~�e��"���,uk�t��US�2�B���14n�W.�:[����ÊXF����6�
�c�>Vy�gX�|�(dB�C�l�z粰À~��^��w�l�vUh�p\0������h���\�g���e�Uq)0n�L�M>���pM�E�h:�8��aI亵ѭ��T|۔]�Fܫ���~��Li^��2I��-w� A�(��?n[�r�-�i�W�����J	kAV�%YK���=}�^w�'� k�D�f��Ժ�nc<�"]�{��7�������݄�.d!�B�#pDGRq�٦�#��c��/s�̯u�°y� A	�:E������l�p�x^5��x�w-�&Zm5�9��ӊ�t-:�9��{�̦�*��������jP{ۜR�A&�j;
nS3����K+:��cV�DO| r=�E���^S�ƇR�	h��9��r'H�<Π�]�T�oY���sl�����Z���V>}V��< �I��Y5�)h
�쎚��tzMl��!�'cJ�J.=�ӨJb�8h�z'x�ၲȾ|�x��\��� �����q�����v��s��+KM��]���&���c����9U��1oB�XN�&0�<���7$D�}��z��/�afC�aa���i������s\"3�Y*�K���A0+��-�WHb�L;]%���� #^���P�)����t��5�F���s9�0U�CRk� �G�O��]�(,���&omS�v��P��63�!4V���
C�*T"���x��`�OY��IlE^C�"3%��N�.`:ǃ�'_���~zŎy�5�ZN�2��4{9|��w-�L��p�Y���'��I�2Ϻ�I��F7�V�数��2(�%����,���9J�If�b�2�	��������3�b	�5<��PX7��H/��E
���A���,�
*
݇_��[���'N����Ѩ>�l����W�����I��(���}������i�"��n�	�w�T_�.�M������*V]B��@܀�����8� ������JW�Uӄ�V�������z�!	��m����^ƌ�5��?r_���ysS�H�GW��ÄRk�nz�o�J�5�=	�}��ߓ� &�/ Z��Ao��,��� 7}/����xSZ���mi5B�O+�ͱO١��m݀'!�6���'闅��c����I;W{���.�i�`?�9�b��R�����DaP��F��Ω̫[9��3yZ���X9��
��@���o��%��5����B���b"�!G'�M��d�,�!�z����z����"H��\���*Br�+UHZ�.̚x����y�`���v�s�z0�"�{4uhJk�n'�+Nsd�y�e����~��n&�1~�<&��r�Zx^��1�Ű�cA�/$�Q��ֳ\g���(��[�p��]���vbٹu`���9��c�Y[�t�4�ܜ<E"NY3oz=��Ơ��cW�0��J����""��	i���K��e��%�	N�6RX0����<)�e���Vq�(ߘ]���MU{�ӌ�&�ۯ����\j��Aʮ�s����*������,�"�V���B��e��P�p!�0S�mf�WXǿ���e����4��A&�a��8�k�0�����@��t�$H���۔�-�A�.�{7~&��h�h%���>��P>�R�z
�֨m̔��d�=��y��+���>���3�?z�Y�fD��)��<�S�#ӛ��C��]�ȍ8	J��n:�*)�r��9)a?�A�� �׫C�"y�{?5��Q��B6/��u�X#a�Ù:߰T��yδP��dq��K�ف�F�{�Jo����z���M���4�'�L�������]�������З�l�FV�IY^$U������������&��;�W(��zdJ��}�:.[�T��R��)�U��_��9k�|Wܥ�tD�N�C���]?���(��=
v���`]mĂ(�5Tw��֊�w)���,�]�m1k�8
2~��1{�)��Q*?��TSV���Ý��C26�z�����Y��w�U�*�$c]��Q7z��|�o�Ո/�U��Gn������*�q�l�)�򡸲<�L�6�D��}�5`!{ɸ/gˡOo�Խ)�T5`��pr��.< > ���Y?��\n|S�{�p�\c!V�Gy��w&�V{��Y��T�(Po��霩�C ̪!�}��o$v�L�e�N�xkf�d� ^�����5���٪��0:����W�h�����GqY<%��\\!l맯�E5��[ @�L@ޚ��P�J�P2 ��<��^���>�.�`'	w��j#��WY�������Z��_[�  �w��
)SD�jf�A7/�;Qnމ�"2���*-����d�ѫ��������Į�87(�DR�����ym�mӈ���gے�!�YH)��l!�b�z���颅p/�8���P�q�:c�&����є=c`>A<D��0n�Ѻ$��M�)luũ�#z�Zr�	Id/|P��������X�qifz�(-W�m1��臫�$�G�~����A�;��Se�����%H��&Y��e?�t|u�x��P�H�<S�_A��J>���w�'y��`�����0P2�p�&�q67d�ۓ�ϧ��C[�U���X���v=,��ySr��~"���*ˎV������0VQDK8r*�~�:qȓQ����?�(����R���X����-�	ο�Á͈dI�J&��x��OΠ�����`I�p��E�m��|�D%oS�P�l[x�GШ`���$Ef�\'���Rhq�)�~Tb���J��?���-���]o�~m'�#��T��!��V�?�עs�����ƠXw��Q�Ek�[(׍;(��B��i�A/����b�_o��t�,�!��#�İ������Qï4O���(cX����ZB�嬩�����y��x�#{��Qpk�D��"��}�QX!l�'�6���c\{�X`�� q]Ҩ�x��gA��#�TѢu�a������p�B�I-	EC��?��!�(��l�s�=����8~�[�B~�yM�)kU59Y��.���QͶ���wX�oE�#V˃͓�R֊��JR�<�VL�ZD_�z�ﲜ����e&9�.n"l}��<Ba�Sc�1Q=M��-�e�fW��o�/R(Yʧ�c>�|��x�q'V�}G��티Wa"��� ��	�_0�I8\�1��Z�z"w�c�>�av�+
��H��)�GE��^VX	�h{5?�	�%t����Y_&�:�wke�Y�Nt�>���gB�X�e�����!���{����0H
Weۤ�@G�PԼ�<�R��k���~�. �)�<Z��Ȉ������t�1�%���=��%�O��T���۔4�e3�����0�|� {�����y����	6��N��w�˟����Z̜���1_upڶx� ��G�pe�w�s_�(7�ʬB��$8Ĵ��KБ�F�5���=���Z���%&��s�����*�b�0��b˷�	d"���b? �G ��(�p���)4�UE�57�V�{����~N�;UmMy�v�O"�m�۵t��]�e�m"i��L%�힉��AБ���q5V�W��	<��A����Bk���O�3�蝥��:vՑ��0s�r��C?CS���>@�7�����-¸�3�M��	F:���ת&lK}u��Y��>��)�E�j�($*��_.�yq�͓�Zn�M�D�]��y���h���U��@#c���oQj 
�>u���C�)���
��y�-��7�&�A�C{�ck?pl�"=_q�ct���4N#�Z!�[K�>l����J��Ғ���M��M�n�o����ǯ��� E��U5�"Z�=�z	�g���C�ڹF�[t@Ƽ>͌�ӟ�p�Вy�p�}+�D��"��".v[�J/�2�I�"iC//j?�6�H���XP��q$�NE�$�]�$.�4�S0��K��b���l�Nj �\���a��H��;)�o�$�>'��^�̧�-�T��k�ۜ�s�/M[=0$��u��<���NOGc���/x��S� X�0|޲�ޙϿ��dM
��6L�zQ�Q��t��4S�G3���eE��s�`н�8�q���҈�3�a���M�B�%vruƚ?XAHS�W��a0ѻY����*�sp)�|�4���Ų�9�'�t{u�}2�߀���/���q�{�9��KcLI�r�����f�47o�q/����@�ϟ"����㱚�h�8B �lK�C��\k���bs�.ڮ�rWd���%�@rp4B�ppom����d�w�yS�A��;	��zP.iuA5G^�����A{��2��C���g5�uک�И'����i��B/�@����mp¦�+�:���dn����^/��SΥ�I�>�r��[�֘�N|�O��������%��kJ��,G�Pz��f��ᗨۂ����oi#���/z�<�W�l>�[$�f�3�|/�YO�S�V.��[c#ӄ�ps�;�-�Q�.y/�;<ȕ�׀ a�"%~ڊ�t�ư̂�r"��:)Z��VI2F�g�Blw.��T4����,e.�B�D�L��H3M{p&`���B�8ٛj�U�|��=1����܈?�o�4�׽D�k��뻚�
0���U?�|�,��'JTм��﵊±[���0q��n]��/�a�����Dɂ�'s���4m��y�O2�)ٍ�>L\�K�����b�Y��In��j��S�[Q2K/X�G�n��r�D�o�0������1�v4�m�ɏ�s��W��zl߲�SE�5K�m�?זQ9�1���au(�����V6���jC�#���f�Zt�]r�f�%ׯ��5��/2ׯ�靗����|�"���l:��E�em��u�O���8��Z
����:ς�u���̷�;�D�U��#+���%���E���.��I	�������"8�u��_ȥSU0�U�@D+BL��#TI�'`��}�ZVҖ���@7N���g�~�����UCS �l��Z>x��i>�֋;"���,�x'ICvֻ�<I�
�)?��7�1b���-��q2�p�r1#%l�T
d`AEp*A�N��&�h�֯ů��f��|��1ap��������2'�{����H��O���
�v�u�ϐ�(G�?E���� �����E��pl���H|�X1	�M���2`�օ&�!Z�:za��?rH����F���b=�������<�+0�ާ�_�����w��$O}��=��}ztϷ�]�떡��Yx�Vj�^��
�.��fs�l�^�k�q���kɯ`�DAh�f�V�!�5�Y�%R����1�sˈl����k�̾�1��w����Qϖ��ss��F�tA���$�bYa��U�ot~16��a����M�7p��A�����*GQUD���6�Z����&ػ�ڦ{j��/�
�M*u$6*�#�g�}M�����/_L��|���#�ܹ�G)'�$�F� �k���=RGH%d+Vv	c���,�Ug�Yv{���QW8�B���(�-�GV0C�[Ǽ�
È	�Ro�ن��A�*����?��.ݏɝ��Q���@3�:9h�zCI(����kױ�sޛ�_��SxDg�������Ky�J�,}��c)̴��x+̚G��s'e�uD|`2'W��Z?G�d����b� �,{e��w����x�K.����3���(���W2��7�LF+�Y&z�@s!�=�Y������Ynк�%�������I�uB��t1�4æM��m��Q�&)'
�q	�4��{��5�%7��[�Ғ1����z��H�S�{M��lD�r�F*����k
n��\�խ��ZewR���Ƽ��͈
������57(��ksv�I�"y��=�	��i�RNrrn�_R8{v]d��9Y�XFQ���T6�_Xd"G�yΘ�Ġ�+� sg���1<���+��|��Nî:2,�l�N.Ћ�>����r�@fr�zwvT�I�.�)��*w���(� ���P1S\�av���/�IQ��:�MH2\^fe�y!J]�"��F�Bl�$[k�x�#�A\'�r��w��$H^�<Ǎ"?o�Q���bqi �n��K��h�f�"��8�F�0Nz�-�QL����$������4]�i#+�eb��r+V�0=D|�]�:��1���V�6U��f��{�qId��ʲ/�U#�����0��uo\:cI)v��ĽG�d�K� 1c�m� �+��FuQ��L{���z��r�CT��6�X^�jp6�ݳ��O�vB���sGR�	�/=@�?�]����r�pKIևM����;�`p�9*1~��ک���e2�0,N�<��|����
����O�x����-&�LT�!��z;�*0Pi���R��$�F��V�� ,������`����n�cj��0!�������1�����&�g`�If~�t�Ni��}�[TĕJR>7���]l ���x��bw=� �;�޳�\�?�vӝ�h���JY�u�
�>��RSO��h΍�D�l�Ȑ�#�<`�vJ&V
�O�b����.~��ݒd�����K��a#��6�6s�Ks�9�F8�>A^J��!h��9@�`�id��)��t�-j��X��> Gܼ~I�6bXp�<$�$WYT���}�|6!y��H�yZ��U3U�iB,�(!�.
�2�����3׌�T���@�wn51���-��,��u��;��'�PJ�˙�����J��P\(�ΰ�Vv ��M�cc1��ԇP�����������z,qAD�~�}��7��O�0.��^S���l���Z���ޏ���8tQ����񣌙D.My��8#-�T��h��[0��ɿ��M�}���i����x��]*�-������="C��*��q���\mQ�u�|o&
u���,�9����	�Af�`.�~{'��cK�f���XL)R��I�b�~|��L+�V��l��{=D�2cI.�U���X#�˞��{�θM�$��Rd��co�_��� v��q��%��m�G!���<�l�&!�FR�z+v�R	,ٮ^Qmc�6�	P~,��U];�A�xW�ǒ�"JR��5ok1��W��U�����ɘ��⨫�t����63��Gr]R0����`���5Ȁ�����2����`v�E�#�B{�!4�>&s���4�tH}�t⺓���M"ˢ"�6��F���6?[�=[�۫%tLa�����V�\�3����I�:0g�]���%��:O��_ n~<�iH��/����mG��Ɏ.:��3���@5O{�ܸ��j"����0A���$���	���~G3�?4׳��6�^vRy�J��%Vh�*\���k�Z")$��d�"$��������\��R�w��B��g�L �J�XB�"���m�΋Z��j��Ɏ���R�������>Fn� v�d#� t����	kn�������-+�V��&=S�J&��N�#�'
��.���R�KMej��W}bYCD��[R�{'jV�N��Bd��fJI_����}QS��*\
���Q��۵6G}�g�%	���[�ciP=�li�#�Bz,�S��l�+嫳��ײ�٩x}w�T8Sw��Iߗɩ��s�W��e��h��A�ǊlT��}e��+[.���og�ue�pG�xQ����Sl,�*�����m?,X��z�p�8Q�l/�>��4�+zA�n��gT�!���â��6��8���3Yѽ�Ȥ,�]�&2�����	`|��8���oW'�����1��^�\�_0O����v�|�7
)�8�U�<�[�6����Xol��F��Y���g�z�fu�ii"SC2ו��G��sE��6"B��q4Ԯ�
GV"�%����ŊĄJ�M��_�� ��S���JVH�n�4ɔT_1�f-����(�Z;�����Kb�G���;�Y�g|"�*X17�g�� t��I�|x�������} j�4'y���$kn�~e��Б��� 7�)8h#G�u�t�_�� ���J#*qe��R��Ȕ|��R����=A�<�`�7'H�)!��d/�mY�A4m�ׇ$/���2�Ӄ* 0����Κ2��6�����J�i���=�1\�q�A	��Ҿ=E	�����⥨smW��%7��-DD��)�k�?�ܶL^��0`:y�Q�Bp*4yhY~1�L5����fs���8���D}$cl|������&L]C�Ң����#�*h:Ԃ%P�r'������:�I!AA��p�I�9��DT��T�)d��O��ujR��t+�6��̬���]1�+��r	�ڔa���ͽ���8�)�Dـ���i�}8A`��s� NX��.Ma���]�G��T��IL��s�ށ<>�CsZ!�l�#_�S��kJ�1�
H��GRyA%�`�������+�j�� ����$��mç�����<�R3O�C2$A�LL�f���.b������
EB�<�&5��*����k�3�}��۷UB�UE�yY��k�b�i��� ��~�2�E��F],���C���D�|�Y�E>N�������#��;��\F��~W�T��tٱLd�IT�#�����	�g�����O����G7���Չ6�}-��L�b7�����T���x��F;�@X�B��G+���\Ţ�":�e+�V�x(�x����E�6�v���{�?�(�E�爅�ɿ���x�x� ߻G
��}�:"4-�h_���7��]��	~���>V:b���bk����F��&핆�J�#�s"ۀʓ��2.�Nw�	㛊L|p�^�W��|���t�@X�.|��BFa�ꚏ.ɘo�Z��g��������S5�.K����A;�K����恬������\�6�di����I�9�=�\�Yyp_�,�gMfn�ĵ�wnҿ�+�}\��74�]O� �!ԱR"���}R�uؓΌ��$t�G�fc@�q�ѨjR��|
���DX��X�4U9��c��ç�!��
�8p��]�n6� I �yeq�O�����$>���:��)^M��������5�0X����j_ �8���������������M%e?1��j�G��RN�Xm�"�k���`�bUt����W��*�7�z~�0�e����1 ���FԎYai��Я�6<W�ٕb=�c���=�TC��s柩��ќQ��>�B�b�P��{'�q�
�;�oҟ�>GRn��'�?o�M~���zg�8�X��'ۙ��՞)m�y�&��A��>4�F�P��m�o	JSh����^���s-\\��c�g1���+S��]�UT��ߙFڅ�]�ty��fW7 ��a.�/�5b#���D���RA�º��*7QC����_x׳�dq� 1>�Z(����l�iu� (�r��1(;�{q���-�Aj
�Q���M���V��	�-���or��)�`dh�/��4c��5D/U��By����/^5�����2Q�4e��g|���,���1���cj�=��c2�_�=Q���r��i��p�T���\�¢�&�7�N�b}�@�.�7;�_������k}sT����tD�&B��� c����52{�J,�&-���p��<wR�;�"�T�J^cuĦ���W0,�Y�2�Q���ԃ�MG7;����C*��cYC���Zo�߃;~z!j�����2��'�w����X��t����y:+l�����a�d.�[z}u�En-Ztt��4$��q�ӻ�t'pMBd�J���
����e�*Y�w�s(ҸY��M�N*.�_!�&��Q�e̿9L{��Tu� �L�X�^n�X�
��.C�P��Y�sdknM��.��g�E�<��aq�X��g���h��h�E20��Q�Ў�T�&90���	?�b�=�|�-�*u0MJV]_�n5�JMu�:�����i��G���M텨u�˅�_�*�c����G
�\x�$$�g�v5��ٻ�ү�yY�J��Jrf&��dOE�wC��,�3�g�$���|&*�8Y�FjSU�s���i��-k�v0��$�1��cT��UeVr�Tӿ:AO����ʼ�wP����j�ݧ��|`�1���P��[A�Ufnm�u2�S��v�����#� ���"6�ٕHb4�0���ȱ�j6�	JGA)CAg��s�i��q-�,�=��{��BHJ�І��%S�a��%\�V����j�tm1C�@���NsyLc��g@Y��&������G�%r�[���j4O7�+�pkI��0��j<��!�O�G.PA���N���Q��zd�̰W��ءu�I����]fSt�8�AS�0A�^��啱�����K����ώCQ�U�3_�<�uf:0W��6˃M��?*�Pm�^��?#}�f��ܯ�W���z=��]M�Fo�!�	�#C�p�T�wd�?#[��#�[چD�J��הfjFs�b��9t^�,8JSP�Oe�2e�M��a��.}��}��U��} ٩��y�Ya�*Gtc+9��hk��\,�/J�S���5#oN7Վ�y(�X������팇Sҙ����z��1�>3a���ٙM\�,4�\�J��P�E�	X�4ή4�W���<ϟ�b#Nu��V��iS��h��A?4\6A<Ό��SDw�h�ґ>��z��ww�D��f^6Dy��Ku��-s��ϨW�����!�xˌQ~��4%:2f3�� ��˲v��*��C㪱ӳ�wR�R,,��bT��ŞQ��XY|a�����h�R{���2����S��m� �lJ�7��[���*�}E��7������P�U?�Y��ϧ_�㣖�v�)��n��y���rd��UߏC�����`�O���Z8�&�(`y�{��h|�ol3����fp� �ar�}O�����N��}�b�!���
崓n$�����;�W����򺞁ĩ�#<�Z����.�TB�<�]MOZ>�� ��^�P�A���+;�8�_��*J�vU�/�� �lS��˧��C&`Q�k�d��dK����;�]�CǮ(%�	>Ɗ��ʔ��0���U�)�PʵH����]���'�,����-���D���4�Y�}l�W/���������@��5D87�,Ǝž?7NI�� #�Q�$~�⯞Y�˔�����`Q��Ҷ�!Ƅ/��Ѳ��0ӊ�2-B&ꀒ� c�yK$@ݺ�������=,v���T)����"]6�vf��3=���EEZF��L�Ӆa�8@���C��b�,����1�i�4�/�p��tQ=dDAN��T���a�ݣX�"�+�#��7<�
���C��	�,-��s��0!�u&��e�}�qj�V脸1Y��X��a�����ܢ�Q�6��.N'�/���m�G�$����͆����1>-�Fz���h��@	6�)+�'�!'�^PU�>7�1�/�Aҽ���ũ�`�]l���+F%�h���]���ȲQ{����i�B���rvpZ�2��
5�f$zQ��(�����υ�Χ^�?�to��+�$m��@�u�V*��w�7;���p(��A�|IO;��JV�'&�^�"/��Ș#���Z_)�_��)J�
e�O��p�׬g�*k@[���y� g
̉RB}�n�X�Z�ow>�m��� ��q��7:����966}79���ަ�a����Ք&�p4j1�+p<���$-B������ֹd���3TQ�b@��ݔ���a��u��N��H+�mS�Ed�ٙ&�`�Q����Os}��E�}����X��F] &xd�Ǳ(.���������eO������q�^|	t�����p�2k�>�������϶�Q�d��x��)�EZ^�k�XuB��ϛ��X`��GFU�R*1�cu	U味>�ڟ�1֟��+O����DOe�No���;v2dn��R����F=li�#j
G[�m��XO�Id���Xz�V�D-�J�4j��h=�^�^n���8��������vRb�*�{l�?��eV�e���a���o\@��𪸨���,b$�%�S��Åघ�%�Q/���]��J���6z�X���H!��])��Q�g(�]6�КW�e��=ef+�ZA@�k�bj���U�bO4u�q�X�-�Jq�6D)�|��%eZ�J�۬$���ێ{�$oU[�����+�B�����cN�a ��`�|�(�c��+p�����L����dͰ�Z�q$L�]񾈬b9����.r�:\�6�����J��lo>�ͩ?l!��:f0@���sЯ��C)��:���}*$�_��ޖF�9�-� l�A���qZ��G��wO����H�_(�+��^����2@�*n:��~���(��k�~�բ|�-@>�(���b�=���|�ޥ��k���< T[@�a�]��V���u��i�d�ǅ�4vm[�;�����孠y����w�f���`Q����r�d^�f���^tLʇTxȲ������ѻ?�/��;�x@|	��>��(�T�� ��������[ag[�3T���¶��|�;^�z�?[�=�pK�$'I<��M1�kp���1�����ѵ#9�T0��؉g�����ؠw0L�"����q�u�d�A����3��*���Μ����ub�ɖ]�7_� z/Sd��l�Mlbښ=.m�v��\�ݓW�-���~G ��l�rΚPi6M1)U��~F��@�Rn���ޓ\��f}��RY#�z����q�J]᭪F溡5N7�jFf+Ys�I����|�p��6��5�;/��&����e7RM���^a0�L������i}�����=a��H`��i�v����2�����a�i4X��ʿ���ȡKP`�A�)�s��w֘*�u��:��4�`�̖����o�8���yPAa��7\������Co�~G҃d%���s%�(���4�l$d���TYPH	+UoE��f��g#<���G`�����e�1��"&�ҵ���.tpc�w2+�CI��N�����l- @G��ZB
��h�4��´�x�9q����G�8H�S�P����M��t�b�y�gW ��t0O�E������!#P���OW���B��	����wR��.���	_83�u�O9��y&�׫����M�e��Yxhv�=yڰM�0T�o�Y���l��9��Ä3�ħ�GQ	���)+�W."]/�C}=�n�P���$�[6��.�Pl��sZ�)]�/#�!�/fj��y�H듼L�y>�A��Pa;��wU?)��N�F'���b��0n�?�־�pHo-�2�Q?4��=�bi]^�"�O�p��qd�iM��ohkGh!�z&�d�p�����H1i��L�g,�7Qq�_\�%�Z�9��6�_F5�86��b%{�K�\��+H�'<g�,�nl���[͞������?7�	���}�s��B:�фb$��M��c\
�!�δ�dym�n���H����}>i�-j]�[�&�2�t�_�iϱG�v`,7	>5��q�JȐz(E�ؚn|�LQE/�e�U=Lm�tm�����"��|~ Nj	��R���$��)�ټtmf�F�6�ݬ9�=c2ybe�p߄�q[��t�S��e��H��H8(C�Ǌ��b���9N,p�h�N���M1�RE�W���i��m�?L-���SS�s��&����kcR:eb��X����h�g�Փ]nA�Afh����0�l^�8 �4LU�?�xP��q�7*����N�L�6�n7?���N�H'J4������CD?�A�eBϙ~��?7c\c2۪�.p�ݓG�%f�U�=6/��Θ�U�s���
z�0b��1�<;4G�/#�	,���r�!4��i��U����T5�맩�#9�[�� a�e~��8�<?6����9�X�y��4sMDV��T���H҃�l��i�3��F�����a���$됷L��kB�)Wv�V�/����H. ����c��ۋ�Ȟ�^�)��ϩ���|Lo���j�p��D+/��9�`�y�:,� �E_'�׭�9ȟ�	~7�jxJP����a@���+=�%82/�!
[r�z.�n�+"\�u,�%�W<𝟅�Y���]{){?o�f� �y�@�X3ı�,y�`�0jU��ce��B�{Ȯʆ��"����o��Hc���?���؍��P����g�,AB��	�n�lklnJt����0��O�ߖQ�O�(�T�b�@����+���F�����R��!�hE�b«����"^��m���{F�_��s�<A �v;���W˩�BG�t��l-z�(HA���6:�0C��b��ȝ@�QS����p�U�m)v�D,�����*U!��Љ�(�C���k��
	.*|.I��AS@��0��c�Rlgv�8�Җ������X�"Ŋ�cy'�^Z;s���k�=��*�r��2LNM�b�՚�Eؼ�Z�C��a[�L5�4]d=?(ʪuҙ�c*ے~��0X��8<�k|&W��ri���
�h��@���-i��O�@P�z!~w����P�*k�?z����(�j���։��?/�:���=g%�$�u��Y�`��6�/.L�/���v�7A��׶��x,�|B��C�q	������{.e��Z��l���ME���\¡!/��@pf�^S.T�6�T��g�o��8Cv���S�->1�
�3�6��R!9���⻬ts5�ʻ���萲I4ѳv+�d��2�
=�j�N`��j�˲�6B䮆�{���l���\�������a|2(,Jt}��&��$>'�fC&3ܷ�{Ĩ4����k�5n~۠�q�gd���i>s}s&�0�^�sO�N��;����_U�޽�"Q�sˁ+u `�22��-���l9;�dd͡ST�P�8������>�p��-9�9c�Z`7C#ޅ$��W"��2]��k�*�s���dt8

�H��#�~=����6}K?uBx���i�����}O�&.Yn�_/���q���t��Q�����["@��Σ��Ntf�"82f����͑{��\�*�t�\B����~x�sz4+�\a����{j,������:��XP�6�����U����*�ys��H�yvf��%�@
y�9����^�Q�y�$���~���z��'�Sh$��_`_��}p���e��#o�J���|oSuQ1������A����~~rl�!9���hĒ7{�5�#[r3�/��ן[I��=�t�#i�o��50)F��e���MF3O��T�vNp�el?�362�M#hт���1��uT�8�#��Jc�%�=峞�2H��:-�����Ѽ���M%)��m��$Ƀέl�r0�n +ֻ%�ؗ:[9L�J�%@od�_�2>�_*�hVA(��@�X�ҏ"7r�-�I_������|��p��R9U�Zok��ư7^!�E��\�G�4�I,��.;�*��EO��SL�h	� 1�Y����䆛_�����B�"N�aH�~�Ĳgo���R��
�?�������@B�GHn��ȗ8mBHZ��?��ڌE�9b��;�������:&%]�����4f����0=CV��v��u�81�qމ�G���V��GB��@Ru`�s	�'��8��������b�����$��*:�/�%1�ii(,�J��T���\#'�>���O�����7�M1 ň���u���)���$]�����#�nV2�~$����J�-��#Ł��ebw0�P��ˇǒڼ�D��ib�� �,U���V'��!:AY����������9�B�)D$f����)�����+8�^-��%@�}ug��]�t�Q���|Y�XZ"E&��k��K���w�����d�;tN�mЦB���J��Kk�T�D\: *���j�?��j�1�	q�~;3\^v����*�%��XH�%�^%A�V��7GI�]:&�ά�L��#��xU�N���o�2�BP�\��m���Q����o��#d���4:	�RX͚��-u�� jxxk�uٝ��`�[C9�K���$��������V}5�B:.�o�*��7K�s70f�gv�<F���U�0y�m��������a��L؝�%w�C�}yܾŰ�6�G��[��*&�5�+k���<����\�<�,z�i lL/�f3SS4�M=�0h5k7,؅zR?���MCJ��?6S��\iq#[�H��3Y��i�l��pZR�/��6��]1@mN��?�8~�{���YD!"�x�n
�R�s;Q�Ft�:�+(����e���+�ln$������d�%~
�`g�q�j�g����c���w��.�'2.N�֕�\���� 4�хG�ЬD��MhmO����]'ա>�S��+q빬��	�� ���ʣ��?�z����+���f��2Z���d^��%�9��u�X��ʷ)2��n�B��H�Z�z�4�)���Q� �U�v�c`6��H�x�q�,v.߾i����j��U�Xk�~��s�O �s� ��GSX����V6�\��[��ZU������^LBw�"O�\&���~�(�~�Cy�FB�9��
22�
��YV�*�Y
�жp�����2�G���S�A����2���������E9ٝT��e�|mm���B�bu~�t���a���8�vQ��;��`�A�D�2��>{�3i\�8�W���P��&p����YfV���k�N�s��\�.0�_�{w
��.��f���=<��vH�G���7�⤍���I�`�+I6R�"D����)}�P���0��EV{���#}�����k����M�����%g�~XB�yo����}Cz"�����!�r2&JUN��44�{B��}���TY��WOE.�L��)l]׷`���`�>U#�i�:wV�MʷQ��2�ߵ���Y*?o�)o\�\9X)�E�3�G�o���D#G���X�-�/�I��j��3k6���Wq�\T�WM��+�ksE+LTG���I>C���tԁ�񋶢q�G/w��g���tK:׏K�n؄N���w]W�[���9T�[,WO�_|1Z��`.n;���c͙Rg��[��(�蛅 �C�MOn[Ob���x{L5��*X�뢔���&���/�էdZQ
u~*��i�������J-V>���y�����M&� �}�{�2�^�J�+�D�KH�f��Y�?�_�]�p�>��Z�3"���`#�y����Rβbܭ�>zd�c��F4=v�R,,d�Q�q=���xU�v��seVG�| �^m�)Mǿ	��kx\iQ�LE��.��0^�0l�81}�Ü��}�!�F��nή�:���W/�P�X���5���t����Öj������TJ������4���\����p�F��μyJf.I���U}��;&�5��R[�m�g���\��1��?��wM��vI�j���ZDzkxs�i�_b�-�|Fh'�X&��<R3�(� ,(u¾,+I/~b��#B�q��Yp�-�`���k�J��C�0�+�'9�6�VI�7�l 8�䗃��%:�GVC��\3�����ëz[e�Vu�0�d��[�XK�b$�v����O!��K�jY��\S�m�媃k����y�y������hv�"FOp
�]_���T���P�D��-y�&^H�̥`�"�{�Uѩ����c&"��㚏Nﱨ ��V7�X�B b��A�2[J�o�Ϩ�VZf�	�.�a�(�� �tC�x@-�/��*}�_K�|�gw}��jz>(dDT��cT�eoV��Y�����M̚|���պ\�䩱Q6�g�FX3U��o;"�0ƃ��Ĭ`%�h"��j��D�y�_���k���l	�+�%7�q�s�9�¨�տ"V5Hъ`yU�.�x�f���͛q&�x��(�wKF��*�J�!k*�����_�ə����#�ñZ��dP��K�<��	�{V��9���~�}	� ��R��`��ˆ�
�2{��:���Gɰ���0��"0�Uq�/��4G�����l4+O���/@K�-���p.C�r�נ�V)��c�qh�A��G#8u�ŉ&����8N��<��HOC��ݝ��* �̫���'��U�j�<�߃"�3h7��j�"`o���o}�D��];˳����V�çm�yK�u�߅���xOEI�	�^װ�k+�TR��iD�,�q�q��4i�	�;�'��m�j�K�-i��S #S�}�qP>[%D��-�T �lƑ�:��>_�nCs��W�  Hǽ,��������F��Rwbr�(AI�tuĚ�b���:�F�G{u�(M��ӡ���H*E�e��������E�)b��
��2]�����_ƐȔ�FD3�������������yqKM�9��&5P��+��L���k;�p�<��"����7�����.��^�QȀ���Hc��=�X(=_�{\�ۗ�?�fɗ��3�^��_�i�`г�c�AL 1�m�@ÃЙ		�!��d+�:;눡3q�u5t+�A�l(v�ɫN
;��Oj�]}���:lv��Y�B���08�ц"������ZjQ���B�+F(����9���M��x�b�-���$cif�s�6��e�i�.O�O������n��]E������3"N��
���kܨJ�_��Q8�<d�"�j������X,����V�8LCϣ9�4��00�pEv� v�� �(�/
s���l m���NO&��\8dz1����������x��7��� ���l�Y�?�v��5
�>f �h�Ifi��a�`� �P�ܑ�n�hh�*v@�\j���c#]�Ö����8�Y�i��S���FۼI7y{pMts�i��ڌ�8�p��|���R�����[��oםb2�0*�B�Wq��.2�@��G�;��$~Y�BI��g����tO�� O� �����a��¬?u�h<s�Y�Lmw����Pm��Ag�{49V�c`&p_}:ԅ�/�oa�w���^�LUwk:`G3�����dW�����&�_���ʇ4���ɿ��P`O0��_�LrI�͍(���a��lHm��a��S�;�K�4������3s�b�9y���K�^4cܩ(��(�t{� ���v�g���cE�c $�l3].42-6M���֌�������?~	*$D��+w;!��a�wg8F�q:ʫ%^M���/EW2��ڝo�0�����zU���*k0��C���`������o�{��G�g����C��Z�HS��#��:1�����\�F2_��2�6�.�cG����G��`���N�49�Z��%�G�X`-�A�	Iב?�˚���e�W�el^�	6��W�=$��4)���/V���*�{+���u��^ΰ�yCR�����������^�|7y�f�r�5�:J.�<�9b�:ZjHӌy�������L��Z-���8��r�%|��L}{���s��m�~�f�sE�C�CS2=d'ʤh��̖���
�dgA��*81���i�(�
�LǾ���z��4N
O]}�}Ü�dQ!�?\y�J��7tC�YF�FQ��j���::�M9�/��Q�'t�^7�&�+|DH=��rp���]dD����bdL�@5��N��{wd���fL�l���ZU�A_���+�Y�v�ı�+�$C���CS�����y�嚽>�C�V�����hx����%'-�_����k�m �Nq��j@l��4��򞇫3�y��%W�*��~�e�.�Z�p))�Q�����i)�����ʢ�K���A���!�ٝ+`�/�r6�7��+K����~ �a `�*P��{^w�{?Z�H�16�_�_l��4��z�A�#@�f�z|��d͡�^�����kؽv3xmy�{g����9�y�%����Q���R#�(��M))AL[������*k�2�dd���t�l{;y��rK/��L����"~��L����-��R�N�(tG�d��������#8�`�!����]���Xʶ�����j�j�#��x�=t�N���eܧ�����ii�y���>>O9K�ƙBP���]�Y0��Zd��])H�^VYY�s؃{`��Z��YHe0���a�M*�D��6�o�Zu$:�OC�)}�V2���Kb4��O���e�_O?ʫ'���|Yh�Z�!��q�����y4g�u�Xy�m����
��ϗ���A)o`zB�%V6csEm˸�C��VP���\�L�D�Ĳۿd4X_0�O��A��/����*h���Ä^듄˫���΢�\" Х�)��ez��{os�C2�������=^P{�ɮ�Od������X�8�sS#
����İ�C-d�ߜ.eL�A�b^��DH-�c��Ç���T�8�T[D�6'[I؆�ј��*ᛷ/��	;W�.k�EU� ���*�e��!\�~8\+�����n��>����q�Ti���Nб�P0Z�~9�Q=!�s:-O����ў��:�{�i�m�B^Υ��2g���E8c��Щ�O��U*_�>�Xqё�/����l��x�
訿�G�>���n_��G��d�]���f|Cb�}�������N\�~�T����s�����r���r5V�x"B�Φ�?�y��xiF⊦�4�`xS3+?��F2�
xUQ���뜠È�������|���+�I�Z@�Œ��qb3y�&����w�S��n�?��Ɨ)S@>8zDv��=%:V�"�(�4�CMv�T� �(�i@��C�q��/�4S�i�D��ڇ+uP���e۳���*���>b�X�&���e�P@ ��ZvB�)��x�ag0��F>>���6$�C�|�$ӄP�7�MPFWn��~B��2�ʌ1.�X*҆A�OH�4&�(���Ч����#�PW��Q��zx�݃���	��ybtJ�CDWw�� Ⱥ:�:|Uu�Պ�L�w�qEu�$(��;�]�Y�U@��T���{�_84�B3N)��3W"�G�>Y��Fh�_�CH/��-�%)�C�1tg��3��ż��$v��בۅ?��?�����c�3�B�w�q�K�ʥV�G��~�id�N ��F���X�jTQ(p�SJ��aN\e�GuU�`�廓���DΧ~T��ہrT��bx]M�Q�J�a�@@����ҫ}��a��t�G�������8�'�VcÞ�S ��'	ep�C�a��U�^����E>��ٻ\c���K����0}�WոN&��]'h�l�./��0U<r��UZگ:����Ó%�9�װ�'p��8�;��WΈ�m��ث�I��D��j�����E�$̪'�[NE�K�� +���i�X�7��<�ރ�E����G��Y�8l.���N�h�L������,�%Z��(�Z^���9�hU$APf�\"�,��Qf����?$�T�N�_Y�ypU����#ʚM�3���C/8�A �������o�_B��~~l��i���Á��7R>?=�hԮ�}�����q����i����4'�qa��iOyz�����Ў�Ұ%X��T��Ü���ݟ���T��zȈ.�V(���U�s�&
Ae�>|�\����Ǵ��QL�if�� 0ԩIm�����͊����3@�F �-GK=�����>���4�^0�/�/�\�+�I����>��*a8�9��֔����^�3C q��	�s�+,�0N����K��S�L�q�3^������p e�6���jA�5qb��ȧ7r�� �MnUkoH�݉�Cm�\O���;]�T1�ξ��G��g��V0���pu�-Y�H��E�{
�e@����O��xhd2�-�"v�o<���ފ�qm��G���Ԋs,��b�)�d6���	�JN�RD9Nw��������}4�lgǋ�ޝm�1Wo�L8�c�uap��8�m\���*�g���yH�p��t��Sa����\u��*}�_Z;��i0�X�<a����֊3uJi��}*���#�����{�1I)�<�Wwe�G���{P�l�F��άHO^����6����-��c����GEi=��uu/��Hl}r��8r�,�]�X�EY?���b�}�a�p�v���� �,�wHl��Ԉ��B[a�;���'��ͭ�0ΕN�"=�BD��h��,-���&��L-p	�HIU.[G��xE�=���.]<������&f�|�6#϶���h.�)Z�����Q{�7ŞC(�a�Q�*j�X7�d�W2�5.;��а��j��
�����ǂ��BR��4�m!�K��]� ��	�^�ȭ��������E���a(ҋ1�(�>`�����U4��Z�ۍ>ͨ���{�QgaU�da9m�V�>Eb�8>5aYTw����d}�a�>�D:T]b�&N &�K���ư�M���t����?�������X�t���Ip>�"_�3�G�+�Cq�CHQm��PP�l�R�2��o\�������PCB�P����������C}f����	��E�l:�2+�6�F��U�`������:����>�'�s�۩ҽSg�s��x˥2!�#�����q��� ת����N����aY�,8؈�#c���W�_h��Z��H_E�� �)_H���T5'ͻEGM��Yp��7'�Dq�=���{(��9��Y����r�"�d`XG�(S(�f��f�7[���rv_�.���^�S϶��۩��5�[��@��Y����d��=Aֺ�S��1�;&���(��'p~��DKAGDpΚY���M�U}p�mD
�G�a�S ��������GL#�.9~�S���F���m�?R��λo�%�P��#��	����U�8�5�@5�U{_�*�_��ND��0����>��X�h�"D�԰�*��� �7tĠ�ݴ�M�̆ѺєX���D�,KyxK����*L Af�������^�i���Yj�3�V�2��Gmcm�����+����:��zN�t�-0�����Pk|?�~ڛ��s�c�4s��� [Df����]dг�0K��Tv��[D���$�A2iMӂ0�3 ^�T0��gRM���/P�m>�
:���>1��wX�n3?·yu'<uk#���F�t���`������R��+߫gs55� �~�s��پ���D�|�;�_��@�xї��0+�R�"�DggX�{�:��J3x�H;�C�\�������<c�}���XK�����vb��oW{N.���k�V�7j�~{|����ۥ���.�Z�@" +*��Ӯ���t�]��0������J�����"Q��7��
F��tm.�TDU�
��2�ʢ���K�@��=)H��w3Ō���R�D��m��3��0
L�[�B<͆�.��@��'a]��b���^z�l��-���- S��H9`�����ӬA��$�)��ie�.&S��g��5W��)��q�φx��C0�|�M�s #���a��L4!j�\�O���h��3Ab�f�Ȇ���
�{�������w��-���
�wd���(|c"j3�A4�[�9�?J�L���~"��4)W8-6���T����M~�D8b�h��1�اw��ƛv!(�EY�-����Vs�����a�r�{rչܦ��[>6�I��2S���7��s(�͉Q7�ٓo��C}���/�A&�lؚ��l��W*:�z���J�����K�ܥ�J�2߳��8x��k�Z �6Z�r^+�YS�����8��J`@Nw�lV�uk��)	�B�;/�w�-���4��G��	l��3�a��A��3���8� 0�ꇔ_��_��{�"[0>_0���zѝ��5L-�2�ӖO��Kr~%=_�2�zͦE�����%�@�Lt�&��3H<.vY
�v�"I�JZ�ޥq�j�2�Y.���d^i=#Q*�x0�����'��������PSf@VҺ��M!5������u	^���&��A��`|��%(\lv��* a������i�ד{�0���
f�[��$�?r��+W��$��"�1)3jVT��}�b�Z�����B�p��Lƿ��eEm��97�gxT� ��?<�vFf@��5� &T�'��R�۬���#�뾓�;h�@�T\y�h]û�ǰ�X#T�"�/)S������J��L�laG,mKu/��j�����7�s��e�'�͸�_Xs�!�֛�e}�t�rY�v�s��.��ȡ�]l��/��G��ś�ب�}K/��4�4����;:;�|*�Jby���}��R��^>Ҍ(�Xd��Si�޿��f�s+&�%�GwS��$�n��K:�]w4�E++s�;���%�5�����rF�z)�4k�F�z���QZ���2z�q�H���WCK���	�zI^1\/�᧔]*��=ɫYB*���"*$rw�0����A���_�b��ǭ.nIG�솶0�?'
}mm�`��;��6����|̷)I���&�G�Pa�n�;�4����w	)&���ӗ���R�7EY���8G��id�?�U�L#U��*�)B2LX,�xIF�eg&�F�
a�5_��_�]�´gD�񋖵-�H�<��!��E���ݎ�
��|���eFk�}��IG>#@��x�8�?\��7J�_�$�5��m)ۣ:BSѪ7�n��#Ѓ���B)D�g��b��h2$� �<{�*�G��w��d���fr����z��4�	ڏ�-�6�"U[#5~ԃ?�~G�<�]M� ;�`ĳ�d��܄zC P��E�\l%I#�Ѻv�3~��3�.5.sK�_OI"�I�x�$%ۭ��D�9v��T���%����ۂ�z�-D��R��˜(s���U����������qW��Y��(�k���iQ(f�U����3�<j̝M�T�+6�UC����J8�p� i�菐����L��=�E�Lk�I�ƞ>���+�5I�����ʺ�M�B�0���]�d'�m"5{�5ܼB�4�",i1"Eύ�*$�|m��y���\��}"�v+�9���e�m�4���TNm�T 9bT�gQ��r��@O�"0I��}wa;��XL��Yq�ڥ�������X�V��Y	ZC�g�ay��~��G w��&_bo�K^G��a���y���s�EQ|�v�C�~7���9���8�(�vRJ�`u��I�y������,1ߔ�!͊��*���V�c���+�M@,��sgp�t|ο{	���t�2��͹�����Q�*�[����#�X������j�������R�p����+���R�-�,���M�ŏ^Q-������R#*p���ʺiO>א��ae̐n�&�!om�&��
>�҂G�r��|j������� �g]v���w��B ��ߎs��f{UY��eK�Ø.�YE�q���jŀ|.��1��W�Ȟ!��ou�����+z�A1a� bS~H!r_���:����Th8�&ԙ�	�u6��ݾb�{���E�������Y��̆���w�����bՕ� T7��9���8�	�
�r�?��N��������������e�z�H���Gß��*�
^-ԫ�s�S�D)�Q	�ڦUzOLۘ��^���q�l��E:)�3�j�Z��5�D��K�ˎҾv���V�m&8Yk���M�sq�x嚿i��/|qQKA"$�p9ϭ7�ϸ�ڢg��V�`�'%I�����$�G��EVQ"��LU퐭�V�����(<�V5CMb��]�����'���O�Ml�!%�'l��}P�!_pPN�|�3�G�w�1�5Q��+#ܚT����(%����_+"����ug�̀-�nr�T'��N�:F
�\��b�/m�39�v��ΥWV�7��^�Z���K�@�<�U{e��u��������i�n@�	�?dzn=# �"s.�(Ҹ[h�8m�P@p����3�����uV5� 8�dR�B0����ꕥ�Bu�g��;�?�\i����.���;8�2�Ѕ��C��$R���4�K�Q-a��*�7�I�W���#��s*p�9�M61�a�|�ώ��Ǘ���3�Z���H�G_�y7��;/	 �Ezp�.���r�(����s{��D��R�I�bl<�N���ٲ�t8�������G64�8�$�/q��Ȣ2������W�k�xz].2Im\�+�y�d���=�1U5y8��a�e�v �_�m�˥�_iR�M)�#R�+�vB��nwr�&�����L��7��*����]����Gu;�_@޸���q�$��u�ۓ��U��;�8��*��x[�v�g��0O�;]ɿ'۝��c����Fz�z�i�ጮ~Z��[��yLj�
�SŌco{t_4w�2z�?Ó@H�r��������
BE��X��tWsQe��V4�,�%���tTI��1 ��[O���h���?j�����^%k�aؼ�Ǒ�L]��(�*��rd�]��[+�<t���#ϢT^AP�Τ3�	�x����<���k�����b$���{^��i�Ę�v �>9DO�3�NAh:.w��h��	,��ħ}�gwT��=�Y���j#O+D���ă!A���e".��!�~�23l,�Y������+H�U77p�q�
�Ƽx�=�YC�Q�]�jR�+�7�/D"RNCc��|��WwS�uC�q���?�����=q�a�K�T��[��uj�`,��a��`rmo����>�y������B}�� ����4tZ���q.��7�`�+����H3$�&!��ؾ�a�~��x(���8`UR%�#`{Ǎ�����z��A�����_N2q��K�3^��u��ʸ�H��^��=*0.�st�K����.��u8ذJ81���"��G�D���6'���K��1��rw
��1'f���~���m�8d�������zVMi)�g����o�췰f9;�<����L͹;D5R3p���|���f�i���.ƯWd�"���U��A��<��+*d�hHU�r��d��)�}c@#:�I4E��� UD��Im0'�l��&�%A^����i����.��c8���Ky*To��.��'~z�j#�n��7��o�9���Ң�E����yA�j1P����Zw��'K%�G�t�[%���).(�w(ꕊ|U�X͝�Y`�~��zg@:q����{�v�>�z�/��&���T!lmjFz�-�A8��zF���c����ā�����8Q���\u+ɚsw���G�9)�vq��q��<W�C�(��\�땛�=$`�N���w>.�*��Po ���=Z�M��)?�(<D�� |��c5� Tၠ�B��1�׵���\Ӭ|���d��0[v5 ��!��F�n�PYK%��T��F���B��+�.�oѷ݇��Q/����c�Rt4a7�-(�q���7�_���C|��p��˹(�W	˥#����O`�\+����::���q�/��+��n�9\��@���t� v�:N�w�k��I��Ǫ�y�R�y��C�Y��c:f
j@/��y�
AA��C�S�h��(���yr����6O�:E6l���I#�?a�Gn���l�`�q���i���+5�`����RU��v�-M�-�̵��F�[Mk�S p�1�ڕ?(�&k�d��:uyL�tßkSS��ȵ�k�"�ky�"�� iV4��:v��]s�[��r
%��dh=]l 4E��>�0	r9U�g�f�)z˯�"�H�>u>�A����I8�?/*����h�M��^����_T�{�����=�����7���w�?���ڻ�:�!]㚷�ըé>�(�K����&T<��z�t=Fx��o���$��w���3W�.������ٟ� � �\��;{�ޯ����u�V6���Վ*������ gI$:L�і�T% ����ܱ����$�S�vl�wE���籠9֗8�'D���_-���CW�;�=q' �m
��3�)A�[�;re�����`��sU�Id����k
��5@�[v�Ha�*�n�MQtl+j�"J	�v�|ˊ��V�@�,
�wm�^Y���7ۄL�L}�:"`����R`}f]I�PT�Ji�I�m�ot�4Ձ��ܡ�;��iFLۜ;PvXM(
9^�����c2��}^�x���~w�� �,�`� 䩵���;�I�I\1�3J��"��5,�n�� ���AzA	OoS)�ʴ�~o���aq"pD���k�\��{y[#W��W�&䦤��(w��b
X�'��A;��L�K�z��PL����i*ڑg�[o�H�i�ѨKYEzA־�K�{7��wt8�C�<Y�������qq����vkޓ��(+ ̖a�`a T)Op���t����Y���# S���h�qދޑ� �\�3{��1�5w"H���1nG�8����7�G�W�vY&��$�)r����5����R7Q�FE���LW0��V�8�u��iJ����X˲�^n2j���'�6��Gް������M��E�ʅm��#8h��G4���r<:��8p�$�/�bKg�1B`�g��.
;Y�K,똰�{��?ɨ\j0�4��6�u�7c���ߗ~�Amz�.��L:q�?D�R��>��p����N���`a�җ�o�K���uNU��'��V��d�^�x�d�X+�G���>=�X��q�+�9k_�*��ж�;k�8\��xSa�yT����

��fRA�R��9)p�#���cK,��0��VW�@%儗�=���p�Z�$���d�n��7��_�L,}��k��Xj�!�2���x�(��xWt�_K! �N�2\�t�u؎O��$;o,u��7�Uʝ�?}V��m�06��kߪ|;�q��3>��Ӽ��X��ٓ���|�+�~�;"1�EV���V�U��+!*�C�Y�pG��[�f�QVE��v,5�A�R��ח���F�����4�F���+�*H��p��>���[��d��Q�9���Iv5��G|�?|��e��(���Q�ŢB�+�)&��Q���v�,q,wX�������VOoPH��k��s�t�_��0U ���m��_�ҭ;��dc��C���$?8=���S<�z��N����P�R/��t���>��Í��J���`���[���_9?

���T�̂�8���e�X�	hɗ����dzEY�<�+m��� ]��H��*s8�>Jd?������S\��6��\��P���/���BQ�}&g3u��`sy��Z��J��Q�� edq�B�UG�� u��A��-?<�����60�fÈ��1��۶K����(̢O�e�.tr���z�n´|h.��S(�~�wP+�ы�� ̡r	��8{:�+��'�%G��5*$~���U��i�o�x� anLݭ�
d!FX���{�k�U�Kֆl8�aϬ:��-)�+�5:�����@�[�H|_���9��$M�dc�UB0�j*J�'/kNnn���5�E���� n`Y�p���vӄ"�L, 싴���e�� Y[R<�y��,f�/����5@����& ��Z�Li����j�t����H);��t8�.g��;�NZףI�j��$���֝����w��KzC7���^�X�U����w�,���??�$�p�W�8��������1wB4�{$�y��3g��3���R~��{���j,z��TS�1(��R��Q2��jI
�7���;?Qb���~n=�c	���G:��T$��Bx.�uvÚg�ł<����xjь^���?�q �q�)l�4�p�j&���]�WIgkv�tR,
&��|K��O�/R'��qÒp~������>��i���#���40�(1���4��YP,�o�e-���I��Sg"&������h5�-X<� �2a;�U|D���y&D�� �t%b�NQ��,�c���&�}	����P�O�b=ixc��Jw4�x?~7�ݥ%��:�T�Ɨ�є��c/�n;�&?�)�/F�8��v�K���ӥ�W�Pү�%=�%K��T#��c4H ���B
	\�;� �`������Mθ0��Pd��l��f��-���v�'L�a��9R�S3�RPh��`�^d��LY ���-���y{R=��1+��s��K;���ݜ��ةJl�{&�_�'�T�l�N`�yػDM�N�J`���T�6ż��Ly�p�I=qe�Zd`� ��f)���"����?'�T�Y"W-.�VWB9r&HT���Z�V��"y�ͤM�4[�'7sq���d��O���}ܖ��q�l4;Cl2"n��ȭ:1��Ƽm}Șٞ�m%�v*iip�)���������nlUWA�t: ӞNM�@-v"]�lȑÅ{n�9$�(�P|�C���-����;�Bb��j�S�����>����{ �>��h�Kږ���Z��
����E�Mȁ+�9Q
KQ�U�G�zV6F,�Zė�@B�r9;e�w���Q�����EZ������4j�������N��c'$����E��v�[��&["�W�q�nߢ�Xձ�q��r7�/�ڵ��Kr#b�5bX����k~P@�&��x���sR}z�*U'wWlg���a�L܇{�qb��z���pR6���8��-��̦��G%�כbp�9�!e���߇��Z#�;/�{2QeVBǩ(����
2�Sؙb+�v́���m��Q�:U�}�����D�]ڧo��.�u���#N0� ����Y8�t&&k�F�(gF~��_�⯁�B�[��������X�U n��Q?�day+��%&uZ��3Xf�O_�������T��Ґ.4�Z�yCg�P(�B��9��K����tCw��.k���A��	����4���,�*���Wߞ�O!��7Vp���O܊X�n�q9AJ��0�RN�m��Ԡ�9zy����K~un���-���HB�T�_�R�=����#=������_ӦN����Vj�7�,*��L��E�Q�n1�{k��9Ͻ��� )WB6�4Sa;19F�1k�Y��.ɸ�)
.�����3�p�xo��/$~	���-0���o��UY�yPyq5H&t�´�����Y����E�YB���A�iG��Pz�G�l��.f ����x�c��%��;��7�nx�v�H(b<�����O�u�es����i���%��N�j��~xN8��%@�JL���1������:zԟ@���۾����s��Sdb�ۉQ4�cQ�3e�0�~�<�&�pF��,g^�7�v�^�!^a�����uz~z-��^��3{ר��Z	R���"fX'������~K��A��Y��^,Ӹ�+}�d��i�N��1\G�#����pwOr�{����YiXc���m�J5o�e�}	4�����"��:o�sw�>�.�hԼ�K'�2 �5N�V��qK *(�E�{Z`�57��kmp��:�o�;'��rY����;�9�11�,p'� ��تſ��/b������wyW[�v"��c�G�ީ�e�h<�/�uc�U�[��̑�b�C�E���E<�މHw�G��� DX�8��B�`����z;t>
*�&h�xy�9��q����i���⬐��~L��b���Y��)���'��;�AZ�z��ѢD-|Iq�� �F�C���zKq��{�_�rM?���x�K`j5u�ܨ;j<� ��,�z�\�G��I��֛��`0��6�5t���s/�-�@lY�$�|��b��X��1����WvZ���l�RD���Y��"Ga2
v���X
$��-���d�Cѕx
�I9"��H;��a�����G���T������f��0MT�C�n&�6��� o�NO��������e�Nq�h��#<h���W�8��߰0\���b�"=�~i��hs��/ͫ��ɋ�V�N�ލ5h�#ײ���9x*O���5�	��E�������?1}{��/��6�'��붉�ۚ�������U��;����8D�=�qsno�بP/�2�ޓE�aK�D�+� b?B'��vi���YUf1�>�S1�C�l��o������穜*��W�H,�x��~j$j#vz�Ctz�ɲiq+�\Z��M �KG�"T� ��h���ho�(zVV��u�f��JH\;n�\R��>�^c,�_n|?�uY��g�A�/3]�:�Ȳ����Y&�-=��d@�Co��2���Q!���$4ǥ�R $?��n(A냇��Y��
Ư� ���^���ʛ�7�-b��N�A~$�H2:=���.��(��z�S����+��e��e�����Hx0�k��b��e���Npc�em�#�Q��7"�y���G�0	�v%�)J5��B�u0��>&�s��2�M�KM����?ω�v�;5h���X_-xi  >�^����s�,�$Ք����V&��v7	�/��#n��g��O/�G��t��*;賘�>�pݻ���x�63�k�EX���X���U�o;J��ӳ��!gT]׉��\�r�KjS� �L�V�&_8޲�X���9�{ӏ����c����t0]�j����I�����ZC��7����|H��?c@�L���n�?d��lU�þ銦h��VSs�����J��l���"I��L��X5��M�19 ���^~��:��%3;:p�ި���Yg����H�5��o_u��o+^���u�/c�*q!�;P�s������֕N��� �Տqcdakɀkƽ/��$Tx�AkS
%���Tm�;:F�����( $�~�@Au/�u�#'