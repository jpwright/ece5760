module nodes (restart, clk, audio_out, sw);
	output wire signed [15:0] audio_out;
	input clk, restart;
	input [17:0] sw;


	wire signed[17:0] vwire_0_0;
	reg signed[17:0] vreg_0_0;
	node n0_0(.left(vreg_1_0), .right(vreg_1_0), .up(vreg_0_1), .down(vreg_0_1), .clk(clk), .reset(restart), .resetval(18'b001010001011111010), .value(vwire_0_0), .sw(sw));
	wire signed[17:0] vwire_0_1;
	reg signed[17:0] vreg_0_1;
	node n0_1(.left(vreg_1_1), .right(vreg_1_1), .up(vreg_0_2), .down(vreg_0_0), .clk(clk), .reset(restart), .resetval(18'b000110001011011001), .value(vwire_0_1), .sw(sw));
	wire signed[17:0] vwire_0_2;
	reg signed[17:0] vreg_0_2;
	node n0_2(.left(vreg_1_2), .right(vreg_1_2), .up(vreg_0_3), .down(vreg_0_1), .clk(clk), .reset(restart), .resetval(18'b000001011000001110), .value(vwire_0_2), .sw(sw));
	wire signed[17:0] vwire_0_3;
	reg signed[17:0] vreg_0_3;
	node n0_3(.left(vreg_1_3), .right(vreg_1_3), .up(vreg_0_4), .down(vreg_0_2), .clk(clk), .reset(restart), .resetval(18'b000000000111001111), .value(vwire_0_3), .sw(sw));
	wire signed[17:0] vwire_0_4;
	reg signed[17:0] vreg_0_4;
	node n0_4(.left(vreg_1_4), .right(vreg_1_4), .up(18'b0), .down(vreg_0_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_4), .sw(sw));
	wire signed[17:0] vwire_1_0;
	reg signed[17:0] vreg_1_0;
	node n1_0(.left(vreg_0_0), .right(vreg_2_0), .up(vreg_1_1), .down(vreg_1_1), .clk(clk), .reset(restart), .resetval(18'b000110001011011001), .value(vwire_1_0), .sw(sw));
	wire signed[17:0] vwire_1_1;
	reg signed[17:0] vreg_1_1;
	node n1_1(.left(vreg_0_1), .right(vreg_2_1), .up(vreg_1_2), .down(vreg_1_0), .clk(clk), .reset(restart), .resetval(18'b000011101111110100), .value(vwire_1_1), .sw(sw));
	wire signed[17:0] vwire_1_2;
	reg signed[17:0] vreg_1_2;
	node n1_2(.left(vreg_0_2), .right(vreg_2_2), .up(vreg_1_3), .down(vreg_1_1), .clk(clk), .reset(restart), .resetval(18'b000000110101100001), .value(vwire_1_2), .sw(sw));
	wire signed[17:0] vwire_1_3;
	reg signed[17:0] vreg_1_3;
	node n1_3(.left(vreg_0_3), .right(vreg_2_3), .up(vreg_1_4), .down(vreg_1_2), .clk(clk), .reset(restart), .resetval(18'b000000000100011001), .value(vwire_1_3), .sw(sw));
	wire signed[17:0] vwire_1_4;
	reg signed[17:0] vreg_1_4;
	node n1_4(.left(vreg_0_4), .right(vreg_2_4), .up(18'b0), .down(vreg_1_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_4), .sw(sw));
	wire signed[17:0] vwire_2_0;
	reg signed[17:0] vreg_2_0;
	node n2_0(.left(vreg_1_0), .right(vreg_3_0), .up(vreg_2_1), .down(vreg_2_1), .clk(clk), .reset(restart), .resetval(18'b000001011000001110), .value(vwire_2_0), .sw(sw));
	wire signed[17:0] vwire_2_1;
	reg signed[17:0] vreg_2_1;
	node n2_1(.left(vreg_1_1), .right(vreg_3_1), .up(vreg_2_2), .down(vreg_2_0), .clk(clk), .reset(restart), .resetval(18'b000000110101100001), .value(vwire_2_1), .sw(sw));
	wire signed[17:0] vwire_2_2;
	reg signed[17:0] vreg_2_2;
	node n2_2(.left(vreg_1_2), .right(vreg_3_2), .up(vreg_2_3), .down(vreg_2_1), .clk(clk), .reset(restart), .resetval(18'b000000001011111100), .value(vwire_2_2), .sw(sw));
	wire signed[17:0] vwire_2_3;
	reg signed[17:0] vreg_2_3;
	node n2_3(.left(vreg_1_3), .right(vreg_3_3), .up(vreg_2_4), .down(vreg_2_2), .clk(clk), .reset(restart), .resetval(18'b000000000000111111), .value(vwire_2_3), .sw(sw));
	wire signed[17:0] vwire_2_4;
	reg signed[17:0] vreg_2_4;
	node n2_4(.left(vreg_1_4), .right(vreg_3_4), .up(18'b0), .down(vreg_2_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_4), .sw(sw));
	wire signed[17:0] vwire_3_0;
	reg signed[17:0] vreg_3_0;
	node n3_0(.left(vreg_2_0), .right(vreg_4_0), .up(vreg_3_1), .down(vreg_3_1), .clk(clk), .reset(restart), .resetval(18'b000000000111001111), .value(vwire_3_0), .sw(sw));
	wire signed[17:0] vwire_3_1;
	reg signed[17:0] vreg_3_1;
	node n3_1(.left(vreg_2_1), .right(vreg_4_1), .up(vreg_3_2), .down(vreg_3_0), .clk(clk), .reset(restart), .resetval(18'b000000000100011001), .value(vwire_3_1), .sw(sw));
	wire signed[17:0] vwire_3_2;
	reg signed[17:0] vreg_3_2;
	node n3_2(.left(vreg_2_2), .right(vreg_4_2), .up(vreg_3_3), .down(vreg_3_1), .clk(clk), .reset(restart), .resetval(18'b000000000000111111), .value(vwire_3_2), .sw(sw));
	wire signed[17:0] vwire_3_3;
	reg signed[17:0] vreg_3_3;
	node n3_3(.left(vreg_2_3), .right(vreg_4_3), .up(vreg_3_4), .down(vreg_3_2), .clk(clk), .reset(restart), .resetval(18'b000000000000000000), .value(vwire_3_3), .sw(sw));
	wire signed[17:0] vwire_3_4;
	reg signed[17:0] vreg_3_4;
	node n3_4(.left(vreg_2_4), .right(vreg_4_4), .up(18'b0), .down(vreg_3_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_4), .sw(sw));
	wire signed[17:0] vwire_4_0;
	reg signed[17:0] vreg_4_0;
	node n4_0(.left(vreg_3_0), .right(18'b0), .up(vreg_4_1), .down(vreg_4_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_0), .sw(sw));
	wire signed[17:0] vwire_4_1;
	reg signed[17:0] vreg_4_1;
	node n4_1(.left(vreg_3_1), .right(18'b0), .up(vreg_4_2), .down(vreg_4_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_1), .sw(sw));
	wire signed[17:0] vwire_4_2;
	reg signed[17:0] vreg_4_2;
	node n4_2(.left(vreg_3_2), .right(18'b0), .up(vreg_4_3), .down(vreg_4_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_2), .sw(sw));
	wire signed[17:0] vwire_4_3;
	reg signed[17:0] vreg_4_3;
	node n4_3(.left(vreg_3_3), .right(18'b0), .up(vreg_4_4), .down(vreg_4_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_3), .sw(sw));
	wire signed[17:0] vwire_4_4;
	reg signed[17:0] vreg_4_4;
	node n4_4(.left(vreg_3_4), .right(18'b0), .up(18'b0), .down(vreg_4_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_4), .sw(sw));
	always @ (negedge clk)
	begin
		vreg_0_0 <= vwire_0_0;
		vreg_0_1 <= vwire_0_1;
		vreg_0_2 <= vwire_0_2;
		vreg_0_3 <= vwire_0_3;
		vreg_0_4 <= vwire_0_4;
		vreg_1_0 <= vwire_1_0;
		vreg_1_1 <= vwire_1_1;
		vreg_1_2 <= vwire_1_2;
		vreg_1_3 <= vwire_1_3;
		vreg_1_4 <= vwire_1_4;
		vreg_2_0 <= vwire_2_0;
		vreg_2_1 <= vwire_2_1;
		vreg_2_2 <= vwire_2_2;
		vreg_2_3 <= vwire_2_3;
		vreg_2_4 <= vwire_2_4;
		vreg_3_0 <= vwire_3_0;
		vreg_3_1 <= vwire_3_1;
		vreg_3_2 <= vwire_3_2;
		vreg_3_3 <= vwire_3_3;
		vreg_3_4 <= vwire_3_4;
		vreg_4_0 <= vwire_4_0;
		vreg_4_1 <= vwire_4_1;
		vreg_4_2 <= vwire_4_2;
		vreg_4_3 <= vwire_4_3;
		vreg_4_4 <= vwire_4_4;
	end

	assign audio_out = vwire_0_0[17:2];
endmodule
