module nodes (restart, clk, audio_out, sw);
	output wire signed [15:0] audio_out;
	input clk, restart;
	input [17:0] sw;


	wire signed[17:0] vwire_0_0;
	reg signed[17:0] vreg_0_0;
	node n0_0(.left(vreg_1_0), .right(vreg_1_0), .up(vreg_0_1), .down(vreg_0_1), .clk(clk), .reset(restart), .resetval(18'b001010001011111010), .value(vwire_0_0), .sw(sw));
	wire signed[17:0] vwire_0_1;
	reg signed[17:0] vreg_0_1;
	node n0_1(.left(vreg_1_1), .right(vreg_1_1), .up(vreg_0_2), .down(vreg_0_0), .clk(clk), .reset(restart), .resetval(18'b000110001011011001), .value(vwire_0_1), .sw(sw));
	wire signed[17:0] vwire_0_2;
	reg signed[17:0] vreg_0_2;
	node n0_2(.left(vreg_1_2), .right(vreg_1_2), .up(vreg_0_3), .down(vreg_0_1), .clk(clk), .reset(restart), .resetval(18'b000001011000001110), .value(vwire_0_2), .sw(sw));
	wire signed[17:0] vwire_0_3;
	reg signed[17:0] vreg_0_3;
	node n0_3(.left(vreg_1_3), .right(vreg_1_3), .up(vreg_0_4), .down(vreg_0_2), .clk(clk), .reset(restart), .resetval(18'b000000000111001111), .value(vwire_0_3), .sw(sw));
	wire signed[17:0] vwire_0_4;
	reg signed[17:0] vreg_0_4;
	node n0_4(.left(vreg_1_4), .right(vreg_1_4), .up(vreg_0_5), .down(vreg_0_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_4), .sw(sw));
	wire signed[17:0] vwire_0_5;
	reg signed[17:0] vreg_0_5;
	node n0_5(.left(vreg_1_5), .right(vreg_1_5), .up(vreg_0_6), .down(vreg_0_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_5), .sw(sw));
	wire signed[17:0] vwire_0_6;
	reg signed[17:0] vreg_0_6;
	node n0_6(.left(vreg_1_6), .right(vreg_1_6), .up(vreg_0_7), .down(vreg_0_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_6), .sw(sw));
	wire signed[17:0] vwire_0_7;
	reg signed[17:0] vreg_0_7;
	node n0_7(.left(vreg_1_7), .right(vreg_1_7), .up(18'b0), .down(vreg_0_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_0_7), .sw(sw));
	wire signed[17:0] vwire_1_0;
	reg signed[17:0] vreg_1_0;
	node n1_0(.left(vreg_0_0), .right(vreg_2_0), .up(vreg_1_1), .down(vreg_1_1), .clk(clk), .reset(restart), .resetval(18'b000110001011011001), .value(vwire_1_0), .sw(sw));
	wire signed[17:0] vwire_1_1;
	reg signed[17:0] vreg_1_1;
	node n1_1(.left(vreg_0_1), .right(vreg_2_1), .up(vreg_1_2), .down(vreg_1_0), .clk(clk), .reset(restart), .resetval(18'b000011101111110100), .value(vwire_1_1), .sw(sw));
	wire signed[17:0] vwire_1_2;
	reg signed[17:0] vreg_1_2;
	node n1_2(.left(vreg_0_2), .right(vreg_2_2), .up(vreg_1_3), .down(vreg_1_1), .clk(clk), .reset(restart), .resetval(18'b000000110101100001), .value(vwire_1_2), .sw(sw));
	wire signed[17:0] vwire_1_3;
	reg signed[17:0] vreg_1_3;
	node n1_3(.left(vreg_0_3), .right(vreg_2_3), .up(vreg_1_4), .down(vreg_1_2), .clk(clk), .reset(restart), .resetval(18'b000000000100011001), .value(vwire_1_3), .sw(sw));
	wire signed[17:0] vwire_1_4;
	reg signed[17:0] vreg_1_4;
	node n1_4(.left(vreg_0_4), .right(vreg_2_4), .up(vreg_1_5), .down(vreg_1_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_4), .sw(sw));
	wire signed[17:0] vwire_1_5;
	reg signed[17:0] vreg_1_5;
	node n1_5(.left(vreg_0_5), .right(vreg_2_5), .up(vreg_1_6), .down(vreg_1_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_5), .sw(sw));
	wire signed[17:0] vwire_1_6;
	reg signed[17:0] vreg_1_6;
	node n1_6(.left(vreg_0_6), .right(vreg_2_6), .up(vreg_1_7), .down(vreg_1_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_6), .sw(sw));
	wire signed[17:0] vwire_1_7;
	reg signed[17:0] vreg_1_7;
	node n1_7(.left(vreg_0_7), .right(vreg_2_7), .up(18'b0), .down(vreg_1_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_1_7), .sw(sw));
	wire signed[17:0] vwire_2_0;
	reg signed[17:0] vreg_2_0;
	node n2_0(.left(vreg_1_0), .right(vreg_3_0), .up(vreg_2_1), .down(vreg_2_1), .clk(clk), .reset(restart), .resetval(18'b000001011000001110), .value(vwire_2_0), .sw(sw));
	wire signed[17:0] vwire_2_1;
	reg signed[17:0] vreg_2_1;
	node n2_1(.left(vreg_1_1), .right(vreg_3_1), .up(vreg_2_2), .down(vreg_2_0), .clk(clk), .reset(restart), .resetval(18'b000000110101100001), .value(vwire_2_1), .sw(sw));
	wire signed[17:0] vwire_2_2;
	reg signed[17:0] vreg_2_2;
	node n2_2(.left(vreg_1_2), .right(vreg_3_2), .up(vreg_2_3), .down(vreg_2_1), .clk(clk), .reset(restart), .resetval(18'b000000001011111100), .value(vwire_2_2), .sw(sw));
	wire signed[17:0] vwire_2_3;
	reg signed[17:0] vreg_2_3;
	node n2_3(.left(vreg_1_3), .right(vreg_3_3), .up(vreg_2_4), .down(vreg_2_2), .clk(clk), .reset(restart), .resetval(18'b000000000000111111), .value(vwire_2_3), .sw(sw));
	wire signed[17:0] vwire_2_4;
	reg signed[17:0] vreg_2_4;
	node n2_4(.left(vreg_1_4), .right(vreg_3_4), .up(vreg_2_5), .down(vreg_2_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_4), .sw(sw));
	wire signed[17:0] vwire_2_5;
	reg signed[17:0] vreg_2_5;
	node n2_5(.left(vreg_1_5), .right(vreg_3_5), .up(vreg_2_6), .down(vreg_2_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_5), .sw(sw));
	wire signed[17:0] vwire_2_6;
	reg signed[17:0] vreg_2_6;
	node n2_6(.left(vreg_1_6), .right(vreg_3_6), .up(vreg_2_7), .down(vreg_2_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_6), .sw(sw));
	wire signed[17:0] vwire_2_7;
	reg signed[17:0] vreg_2_7;
	node n2_7(.left(vreg_1_7), .right(vreg_3_7), .up(18'b0), .down(vreg_2_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_2_7), .sw(sw));
	wire signed[17:0] vwire_3_0;
	reg signed[17:0] vreg_3_0;
	node n3_0(.left(vreg_2_0), .right(vreg_4_0), .up(vreg_3_1), .down(vreg_3_1), .clk(clk), .reset(restart), .resetval(18'b000000000111001111), .value(vwire_3_0), .sw(sw));
	wire signed[17:0] vwire_3_1;
	reg signed[17:0] vreg_3_1;
	node n3_1(.left(vreg_2_1), .right(vreg_4_1), .up(vreg_3_2), .down(vreg_3_0), .clk(clk), .reset(restart), .resetval(18'b000000000100011001), .value(vwire_3_1), .sw(sw));
	wire signed[17:0] vwire_3_2;
	reg signed[17:0] vreg_3_2;
	node n3_2(.left(vreg_2_2), .right(vreg_4_2), .up(vreg_3_3), .down(vreg_3_1), .clk(clk), .reset(restart), .resetval(18'b000000000000111111), .value(vwire_3_2), .sw(sw));
	wire signed[17:0] vwire_3_3;
	reg signed[17:0] vreg_3_3;
	node n3_3(.left(vreg_2_3), .right(vreg_4_3), .up(vreg_3_4), .down(vreg_3_2), .clk(clk), .reset(restart), .resetval(18'b000000000000000000), .value(vwire_3_3), .sw(sw));
	wire signed[17:0] vwire_3_4;
	reg signed[17:0] vreg_3_4;
	node n3_4(.left(vreg_2_4), .right(vreg_4_4), .up(vreg_3_5), .down(vreg_3_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_4), .sw(sw));
	wire signed[17:0] vwire_3_5;
	reg signed[17:0] vreg_3_5;
	node n3_5(.left(vreg_2_5), .right(vreg_4_5), .up(vreg_3_6), .down(vreg_3_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_5), .sw(sw));
	wire signed[17:0] vwire_3_6;
	reg signed[17:0] vreg_3_6;
	node n3_6(.left(vreg_2_6), .right(vreg_4_6), .up(vreg_3_7), .down(vreg_3_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_6), .sw(sw));
	wire signed[17:0] vwire_3_7;
	reg signed[17:0] vreg_3_7;
	node n3_7(.left(vreg_2_7), .right(vreg_4_7), .up(18'b0), .down(vreg_3_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_3_7), .sw(sw));
	wire signed[17:0] vwire_4_0;
	reg signed[17:0] vreg_4_0;
	node n4_0(.left(vreg_3_0), .right(vreg_5_0), .up(vreg_4_1), .down(vreg_4_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_0), .sw(sw));
	wire signed[17:0] vwire_4_1;
	reg signed[17:0] vreg_4_1;
	node n4_1(.left(vreg_3_1), .right(vreg_5_1), .up(vreg_4_2), .down(vreg_4_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_1), .sw(sw));
	wire signed[17:0] vwire_4_2;
	reg signed[17:0] vreg_4_2;
	node n4_2(.left(vreg_3_2), .right(vreg_5_2), .up(vreg_4_3), .down(vreg_4_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_2), .sw(sw));
	wire signed[17:0] vwire_4_3;
	reg signed[17:0] vreg_4_3;
	node n4_3(.left(vreg_3_3), .right(vreg_5_3), .up(vreg_4_4), .down(vreg_4_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_3), .sw(sw));
	wire signed[17:0] vwire_4_4;
	reg signed[17:0] vreg_4_4;
	node n4_4(.left(vreg_3_4), .right(vreg_5_4), .up(vreg_4_5), .down(vreg_4_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_4), .sw(sw));
	wire signed[17:0] vwire_4_5;
	reg signed[17:0] vreg_4_5;
	node n4_5(.left(vreg_3_5), .right(vreg_5_5), .up(vreg_4_6), .down(vreg_4_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_5), .sw(sw));
	wire signed[17:0] vwire_4_6;
	reg signed[17:0] vreg_4_6;
	node n4_6(.left(vreg_3_6), .right(vreg_5_6), .up(vreg_4_7), .down(vreg_4_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_6), .sw(sw));
	wire signed[17:0] vwire_4_7;
	reg signed[17:0] vreg_4_7;
	node n4_7(.left(vreg_3_7), .right(vreg_5_7), .up(18'b0), .down(vreg_4_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_4_7), .sw(sw));
	wire signed[17:0] vwire_5_0;
	reg signed[17:0] vreg_5_0;
	node n5_0(.left(vreg_4_0), .right(vreg_6_0), .up(vreg_5_1), .down(vreg_5_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_0), .sw(sw));
	wire signed[17:0] vwire_5_1;
	reg signed[17:0] vreg_5_1;
	node n5_1(.left(vreg_4_1), .right(vreg_6_1), .up(vreg_5_2), .down(vreg_5_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_1), .sw(sw));
	wire signed[17:0] vwire_5_2;
	reg signed[17:0] vreg_5_2;
	node n5_2(.left(vreg_4_2), .right(vreg_6_2), .up(vreg_5_3), .down(vreg_5_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_2), .sw(sw));
	wire signed[17:0] vwire_5_3;
	reg signed[17:0] vreg_5_3;
	node n5_3(.left(vreg_4_3), .right(vreg_6_3), .up(vreg_5_4), .down(vreg_5_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_3), .sw(sw));
	wire signed[17:0] vwire_5_4;
	reg signed[17:0] vreg_5_4;
	node n5_4(.left(vreg_4_4), .right(vreg_6_4), .up(vreg_5_5), .down(vreg_5_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_4), .sw(sw));
	wire signed[17:0] vwire_5_5;
	reg signed[17:0] vreg_5_5;
	node n5_5(.left(vreg_4_5), .right(vreg_6_5), .up(vreg_5_6), .down(vreg_5_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_5), .sw(sw));
	wire signed[17:0] vwire_5_6;
	reg signed[17:0] vreg_5_6;
	node n5_6(.left(vreg_4_6), .right(vreg_6_6), .up(vreg_5_7), .down(vreg_5_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_6), .sw(sw));
	wire signed[17:0] vwire_5_7;
	reg signed[17:0] vreg_5_7;
	node n5_7(.left(vreg_4_7), .right(vreg_6_7), .up(18'b0), .down(vreg_5_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_5_7), .sw(sw));
	wire signed[17:0] vwire_6_0;
	reg signed[17:0] vreg_6_0;
	node n6_0(.left(vreg_5_0), .right(vreg_7_0), .up(vreg_6_1), .down(vreg_6_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_0), .sw(sw));
	wire signed[17:0] vwire_6_1;
	reg signed[17:0] vreg_6_1;
	node n6_1(.left(vreg_5_1), .right(vreg_7_1), .up(vreg_6_2), .down(vreg_6_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_1), .sw(sw));
	wire signed[17:0] vwire_6_2;
	reg signed[17:0] vreg_6_2;
	node n6_2(.left(vreg_5_2), .right(vreg_7_2), .up(vreg_6_3), .down(vreg_6_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_2), .sw(sw));
	wire signed[17:0] vwire_6_3;
	reg signed[17:0] vreg_6_3;
	node n6_3(.left(vreg_5_3), .right(vreg_7_3), .up(vreg_6_4), .down(vreg_6_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_3), .sw(sw));
	wire signed[17:0] vwire_6_4;
	reg signed[17:0] vreg_6_4;
	node n6_4(.left(vreg_5_4), .right(vreg_7_4), .up(vreg_6_5), .down(vreg_6_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_4), .sw(sw));
	wire signed[17:0] vwire_6_5;
	reg signed[17:0] vreg_6_5;
	node n6_5(.left(vreg_5_5), .right(vreg_7_5), .up(vreg_6_6), .down(vreg_6_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_5), .sw(sw));
	wire signed[17:0] vwire_6_6;
	reg signed[17:0] vreg_6_6;
	node n6_6(.left(vreg_5_6), .right(vreg_7_6), .up(vreg_6_7), .down(vreg_6_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_6), .sw(sw));
	wire signed[17:0] vwire_6_7;
	reg signed[17:0] vreg_6_7;
	node n6_7(.left(vreg_5_7), .right(vreg_7_7), .up(18'b0), .down(vreg_6_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_6_7), .sw(sw));
	wire signed[17:0] vwire_7_0;
	reg signed[17:0] vreg_7_0;
	node n7_0(.left(vreg_6_0), .right(18'b0), .up(vreg_7_1), .down(vreg_7_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_0), .sw(sw));
	wire signed[17:0] vwire_7_1;
	reg signed[17:0] vreg_7_1;
	node n7_1(.left(vreg_6_1), .right(18'b0), .up(vreg_7_2), .down(vreg_7_0), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_1), .sw(sw));
	wire signed[17:0] vwire_7_2;
	reg signed[17:0] vreg_7_2;
	node n7_2(.left(vreg_6_2), .right(18'b0), .up(vreg_7_3), .down(vreg_7_1), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_2), .sw(sw));
	wire signed[17:0] vwire_7_3;
	reg signed[17:0] vreg_7_3;
	node n7_3(.left(vreg_6_3), .right(18'b0), .up(vreg_7_4), .down(vreg_7_2), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_3), .sw(sw));
	wire signed[17:0] vwire_7_4;
	reg signed[17:0] vreg_7_4;
	node n7_4(.left(vreg_6_4), .right(18'b0), .up(vreg_7_5), .down(vreg_7_3), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_4), .sw(sw));
	wire signed[17:0] vwire_7_5;
	reg signed[17:0] vreg_7_5;
	node n7_5(.left(vreg_6_5), .right(18'b0), .up(vreg_7_6), .down(vreg_7_4), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_5), .sw(sw));
	wire signed[17:0] vwire_7_6;
	reg signed[17:0] vreg_7_6;
	node n7_6(.left(vreg_6_6), .right(18'b0), .up(vreg_7_7), .down(vreg_7_5), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_6), .sw(sw));
	wire signed[17:0] vwire_7_7;
	reg signed[17:0] vreg_7_7;
	node n7_7(.left(vreg_6_7), .right(18'b0), .up(18'b0), .down(vreg_7_6), .clk(clk), .reset(restart), .resetval(18'b00), .value(vwire_7_7), .sw(sw));
	always @ (negedge clk)
	begin
		vreg_0_0 <= vwire_0_0;
		vreg_0_1 <= vwire_0_1;
		vreg_0_2 <= vwire_0_2;
		vreg_0_3 <= vwire_0_3;
		vreg_0_4 <= vwire_0_4;
		vreg_0_5 <= vwire_0_5;
		vreg_0_6 <= vwire_0_6;
		vreg_0_7 <= vwire_0_7;
		vreg_1_0 <= vwire_1_0;
		vreg_1_1 <= vwire_1_1;
		vreg_1_2 <= vwire_1_2;
		vreg_1_3 <= vwire_1_3;
		vreg_1_4 <= vwire_1_4;
		vreg_1_5 <= vwire_1_5;
		vreg_1_6 <= vwire_1_6;
		vreg_1_7 <= vwire_1_7;
		vreg_2_0 <= vwire_2_0;
		vreg_2_1 <= vwire_2_1;
		vreg_2_2 <= vwire_2_2;
		vreg_2_3 <= vwire_2_3;
		vreg_2_4 <= vwire_2_4;
		vreg_2_5 <= vwire_2_5;
		vreg_2_6 <= vwire_2_6;
		vreg_2_7 <= vwire_2_7;
		vreg_3_0 <= vwire_3_0;
		vreg_3_1 <= vwire_3_1;
		vreg_3_2 <= vwire_3_2;
		vreg_3_3 <= vwire_3_3;
		vreg_3_4 <= vwire_3_4;
		vreg_3_5 <= vwire_3_5;
		vreg_3_6 <= vwire_3_6;
		vreg_3_7 <= vwire_3_7;
		vreg_4_0 <= vwire_4_0;
		vreg_4_1 <= vwire_4_1;
		vreg_4_2 <= vwire_4_2;
		vreg_4_3 <= vwire_4_3;
		vreg_4_4 <= vwire_4_4;
		vreg_4_5 <= vwire_4_5;
		vreg_4_6 <= vwire_4_6;
		vreg_4_7 <= vwire_4_7;
		vreg_5_0 <= vwire_5_0;
		vreg_5_1 <= vwire_5_1;
		vreg_5_2 <= vwire_5_2;
		vreg_5_3 <= vwire_5_3;
		vreg_5_4 <= vwire_5_4;
		vreg_5_5 <= vwire_5_5;
		vreg_5_6 <= vwire_5_6;
		vreg_5_7 <= vwire_5_7;
		vreg_6_0 <= vwire_6_0;
		vreg_6_1 <= vwire_6_1;
		vreg_6_2 <= vwire_6_2;
		vreg_6_3 <= vwire_6_3;
		vreg_6_4 <= vwire_6_4;
		vreg_6_5 <= vwire_6_5;
		vreg_6_6 <= vwire_6_6;
		vreg_6_7 <= vwire_6_7;
		vreg_7_0 <= vwire_7_0;
		vreg_7_1 <= vwire_7_1;
		vreg_7_2 <= vwire_7_2;
		vreg_7_3 <= vwire_7_3;
		vreg_7_4 <= vwire_7_4;
		vreg_7_5 <= vwire_7_5;
		vreg_7_6 <= vwire_7_6;
		vreg_7_7 <= vwire_7_7;
	end

	assign audio_out = vwire_0_0[17:2];
endmodule
