module read_swithces (
	//CA Rule Entered on Switches 7:0
	
);

endmodule